��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3�[�����Pٵ&�����''�qe�-�?
�%w$�W��[��m�w�xH�O�I�	�@����[oVʭM�A��t��B�gx�K���8C��G#h�̾cZ���8���L1�}�L�RZ��L/��W�p���;lB��*�Y��4�%]�Y�:�b�\Yv_f��!P�{
2G�-�Pi���xhB�ё�&���7`��G%����U�^�9���t�M� ���X3���#���u�鉾μr|Wh��h��Kɟ������cG:��9J>:���ϔ"��nE��2�����>pS4s��	�(G4{(S�L�:U�.@�|R0�L8������j��IB�"���N������ys��ė/,ҊN	qh,���2c��-� ��͉��o���a���dsv��s)��.i�}����К0��8õSd A��Љ(�[��#w�eފ)jf9��������-�-��g"Յ}�"ȄP�����}�߃@/�7'�A�9T�)���zG ��k������h���/2A���z�;�-� w���bQ�Ds��?�]���ШM�3�#E�|J�~��'�m��o��0�	 ����� �!m{_�E%�r���]-�O��ΆxI'f�i6�sZ�MJ�{�i�7+�K�:]��u
�qo"�T�wg�õ�6��t��\�K����;9�����X���wH?y-�c�I�{7�|�F�D�ܑ8�g��٧�0�]�� �O>A�\<� R�A�.g�4."�.X�`-��H-F�vw�-�$��l0���ez�U�7�L(%.V���P�S��7.h�ɷ�vʝ̵	W[pP ��[�ʣ�6��V�Ѻ�&�P�Eu��׶��%�\Pi�M7=�h�T-@bm�Q�~֦ I�^�ѹp�	�F���)T%��n�d�r3�H�X�/'���xP�&fʪ��U�(�r	�߈��dkג�Gy�L�6o�2�l���B�	b�4?Ύ[���b{üW� Ī#g�u�Q��H�ޜb>����	I|MW�9�Rv@��Sk`sT���#��P�8L�f�qȇ �򂸾Y1W�I�<���P�|�W��rJ�J�bnU>�G��n�YB��_�5��@�K��s�,ǎ�������$��� ��7 ��A�у�t�v肥�5(ɦ����t�T`�v�WMV��q�Q��f���b����?8�ٟc��T 7�m&]�)�F���YU��Eq�@!�����5צ�^l���es�m_�O�q0�-��g�[A����F{�_m�s)� ؐc�U��	;ݬ���;൉a9w[_ԅ��0J������p�����>�$-op3ڿ����%( �w��׌Og
�~݋�<󹨿���:�	I�z���T�s�r���_�rf~�0}- V�<�/\��'.���L��#�& �KR�e���e$U^�V�KN��� 6�ZX1��� �k��fI@2��)n�Ngː�](wV(�����G��8|���1>�v�=�u?ٱ�v������ʜث������_d��9�Mh*z2VD��:�Ĩb�O��3�^9���<��7�n�(E/�����V�����yX�J�c�h�a���Ph.;��6a-���nz��(��< ��6��)�.�+�g]�)�4<���5�+���{�c	m1��4�Z'V6�U�!�I�s[w���)B�~
��<a��������Lsd�&����BZ�-�T*wƧ�xm��Ǻ��v�T�-$�'vo;��:k+���� ��!�p�[6f��o��L/v� ���!��%*SGư_�` QQo��Eom	��p�J����m]L�r00cwU���(���r�����;Ȋ���P�����$���Z�i���8_-�s4B��n`<V�����!ק�j��7e��#���q� ���R��BU���u
�F� �9��⾤� �[��P��ꣿi��Ŷ�j��)}�n���F;*'�͜L�Sh����e6�>EN���<���$ik���q3����C�5�p��#3Q[��_K�V�;����A`鬳P~�U�����vy��x��W���ȄJ ��Ń7ܮ�#�6�mgΙ�`��Ao�܋�5��,Q&�4�aC��G��:'u{Lʑ�x�E��eV�}�$Dl����q�5��ͮ�a�|(��w���p[d�+� S�,�ѤX�� h\'�_"|,`�숰�(y�著����5g�����;D����`ܴ�P�*�����o�Pd���$/��9n�z�4�M�h�@�6� /ti#?����I���?���w �4cN��b�Y��\�m:תn����'�e�'�鹫/;E~�da�w�h���d!��,]�9�/t�;:���oY�zD��*�����6?m��1�<_���"�N��#�����;�fI��h7��κ�h��P��L bf�����h�.{G'���ԩ���ɮ�㡈-m�Mz񵬤��a���Ɵ���<,�t�y�A�|FSh[�s;<= <�\/��g�(X��u�s�N��DзFﭿ�^�O(k��R2�V@[�'vR*���X���tSp����Ƕ�5�˜�ա3�Jn��8��S(��_N� @X�k����&�^F��"ױx�Y3%�[0�ojG_��6$�x�]�[}�z�2"�k5�q���+����wv5��w�`$�[E6�8�j�s� l�ڿ}���A��*�X�Qe�5�	[�SC�<ג���dЗ�/���]<���q<��'L�B��H�^���~��������"8U��b����w-�
qbhr������j{�(N}���G����Ԑo�0և)6��������x������g���U� ����UNn�AR�Sm�ͶU��?]Ar���"�6��؟�Ճ���v�z���	F���Oj���Z�F��Գ�A��_8��1tf�@�&����[����N`J�g#or��i3��Ha@�ֺIr�M���6�J�Jә���ya�0ͫ�kY�27^?�9٘���A�5a��'�z�Dg ]6N�����k�t����@����K��o*���H��&A��J�$��!�^�<�?�t}��N��
��@P�:��N�.�r�b�y�Z���|]
���|I�y�B��ɐrkj�3<o&7�_3��N�C���C㾿7���\�.���cjf�O,�,�y�i��9���x62�S�ơ���������NCk���#t�v�B��7�jY:���^�2cc"j��:����Ē�wX�� )�aC2�!�9w
Wj�'qy�PAf����J�g�i����t*5�A����|��DC{JE+UO�Yb��l:�0H��H���I���%���3.HD@��B�É�ߕp���۾��7ĉ��*a�&n��D�V�N�5����m�q��c`3�i���H��c2�|i�P������"{ɀ�_*V��>1����)B� :�����xG��S����Se��o�:~s2}�w�5��^�����Ư�N{�}1G����T�A}��Ŧʦ�p�E�5g(���_~~�a�[�
C�
m��E�p;=���#m.ٸ#�<�	�G�S�X�����:ϵP(M�还���di�[��G����NO�>iJl���k��B�qw�O��&c� �����(�O�;�
���5���zިQ
wT��~���[_��(����Aa��1�p���J�t��h~t��\�ߜ�iܯ�o/�(�R�2�\��O�B��ա������<Z5�\޿��O�Hq�~�Oc��ܹ������r������׽g�*҃�(<�l7����Z�����	�m��2O����g.�5�
��~d'�<�y��6����T��cY_��y��?Ī2�<ql�:~i���GS���G�\�bq�["�f�!wj����!�ڗ�iπ���%��U��,l>�v���\��	�dC܊�K��g�)Jw���c����>���������a�jט]@A8�BZ	�z��AE��w7��u�g��
+|�$9d&�z���L��?s���d|�#ϸ\c��vj�ttc�e����^��}Z�g�!�ڀ���*4]6\�8�Z��8Ւ\��r��O��?�g�����/����?2��!YU��3C#�T�O�Ck�HW�Ea*�]�����`6���%S�c׸@}
gOR�v��9x]ƞ7-��cV�����P1,#�Vͣ�����0��i�":"������yo���&�c��my9���Y�O��^/ޭ �
�~XC/�(
�A�;^s=��+R�]��ֱ�N�����>�R��x�?��� ���h �1*[�@-��Ě&�������T_�8�#~}靏�>��B^�����L�';#����1H��Kfo�k\c���,���O�&���[�"�WI�	��]��k];�Q���HE�LHLu-��]V��1w�<?�~��\��5�=K�9Ǝڱo�FЧ���T[�˖�>^�%�Dǘ�j� z۱Բ0��Xɏ.��}~S-�*2y�˶�Z�����Д�4�A�Ɠ���Mt5�(���&y3���]&�����ኙ_�,:����\+�i� ����#9l&P�C� ѡ@��a-�L����{s�j1�I��^���EYp� h�����Yt2����iw3�̂5h��ƞE
�5?j?��)����Óx��i��V�͵0�c/n�6�-��}�R�O�B����;l�6!/d�j���trF�}cZ7)��-�>{h���gj)i})��4$ම���V�ldNq�D�����r��D�x S�����H��:��	�mKѳs�����c<p���X��Sl�#��:`)��o���c�K?&J�R��'|rCLBfi�m��-��v������0�F�V$6��P�|�.z�����}Lr^5)��E����n˼Lk2J���s�9ߘ�7<a�z.aZQ��>�䚸���tҟ�^6�.Sf����5����*���*݌�;��CQ	%�[ڎY"��t��)��]XnWL�����f���<�,M�+�?�C!ަ"t��
�� >�M�U�ž@p�^���wؐoGn�W��(4��yi]g���o��t/%����zp˫_�h%3Ql���9~���ܴ��z\��km5�g=,��I&���MӺ�%
�w7���BOҮ��E�Ё������b
 ��-n̶�	hI�'�O�K�؛�~�-m����+d�[�3JA�g�:�k�gEض�ش���&�a�.�)�'�R�(�޵�P݋:�Д�#�;S�鲞��󑁧4��|�)��1x x�OAN�e�v�Œ$8��ʪ���"bË��@Z��+�n��k�A������y:nO�ND��I*�I� �[�?�K�r�NI~�(��~���N�{�&�P`�XuUG�F��隈�Iz'a���u��+�5�5$Z�Q��	U`�Q
g��6��b����Ũü{ק+�gA/"���D�#R�N��7T��ƶ�6F�+,��f������`8�T(m�=�� S7y� ;�8K:�h��Si눙d:%�OZ;�*���28�p��X2��R�%�wS�eȿ��1)� �a�WUq�C�A{�<��o��Gm:�~��+a	@K���;(iY���7���_z3�����؄|p��UF}��������V���,���ʰ׈�{��?�`�i�HI���V`��+�W+�@�,눠ݫl4b�$�w�H[-�>�X���!��D�Z������/�Aj������dV����3w?���cū���fo^a�xI�����卥�&�)o��N��N����q�r�+Q)�/����U��=$�=�0M����;w�~�h!>�����-9�������̞�C�<̯�S�)��cVY�`r&��4ũ��Ѣ3 A�(O��X���
<����G�gC��*�2CHN!������Ĥ��I��љa�������$�5�K�(i+� �!e��1�K����4�	�����ྏ}z5��c��&��{�`���H��29��2��-���z�������L`���Шl��Lu���~��)��psX���?S�S�r���)��	L"�ψL;�W��8j}��@5���? =��z+����5��� �z����!CF�~`)��.9bw�T:l�%�`u岄-�}��P��:(&��-�Y�M�x=6�%[�=���=ں��Z�%"�����%��?ɾ���C�R��B�A��+�&[ͳ� M�9�B*�Ƀ�+#��L�Y6RU%q
Lr]P�F*ř�@��\�W��_5FN�&�6W�8[�f���pd\�� s`��lBEv���d�!Nb�q�7a�j�f�r�r�����)M�Pdj�KPN�.$�o5�#)�f�r�ѳ6����60�����D;82�S��(�~_����I�ő�-��_t��ų�6m��*�{���ھ^dB��φ;���<�E���`�ktxО˝�����zy���~�n��^T�p{�����~�[�w2��6�3x�P���R�h��j7����'N����2��������N�����ǥc������:�|#U�C�����J���8gѡ#��}eq��*�cU�8C��&�7Ml�[��H0� Śqg�x�*r��$���i�� ȶ���R��n�?ݕ=���1�|ud;@hCAe�ܸ��C.��!�MƩ�����:Tw��3���g���]�rǸ���SEG�6�8nvT�Pc�+�*���%zo&�9a���<_K�S^�����x|���2��s��W`�������g��qvD1C���FW�q��ߒ}3_k&0��(��;�m���f)|�LB<�liq�O�\qaZ`�;.���h��ڳ�xO��� �w\���,ׁ6C"ϙ�I���Ԁ؀aB�@~{����$����Fxx>�yH?:^�ఆm�IPy��+Fz��n�	ڡfYysS[ւ��u�>2ը�K�'�����h�>� ��`�pЃo�{U~7��.�/�g�o�H(�ȹ����7�{���/�c���Z�J��	�&O��V��K����%I{e�W�h��2���!/Ay/x���":�w��;��?5�) @�b'���0˹�^.�R��L�����c��L��$�y`��ߓ���?=��؅T�p�p��+h�҃Yp������?������I�Ϸ>·1�	t�u+�j?I�r2�6P˪3���a�D)�A!�#����J��2kvG�s���%��~�B����,w'-k]�	$�Z�s'��t���]��.E����z{����D��w��n�ܤ}�Q���w�@r0m�����!zwc��,��\ε�aA�W����TT2ȆB��~�T]!���>i������k�e���/���'�s6m{�"��^���ahr/J��|�&��w��
�Pӂ����s���E������Q� ]m�|P�QË�I�� �,rＦhwɖ���e0^��6)Q�|<OK���]��R@�1��D������8�ŗ��z��L2��M����d��	)¢Ә�u�qf�h��D��a?d��9C�< �� �9
���L����T�b���`5��O���p
���X�P!T�2�~�2��K���ۤ"{����q�\�F�phl�����Ԋ�����c��5�gSc�4��������*q�ԅY
2�,V҇���#+g��^��x�X�p$�c�n����W�!C;G��,EN%ԩ������p��f����ju�	�H��fK:��x]�/�@vp���0���f�ii�s�"Cw�N�A#Y��(��|�e@~�X�6��	�I]���{�#1%Tm�3�qm�P��y�֟�w���c����mj`?��W�kG���41�r/"a�1c��ٴ�Y����4C��	F���mӱ#����Ԃ2�Cs&����g�76|�6����[���jN�23o�����C�&� �I�KI��oR�8]�9%��n�bh�T`}3��/N�Y`� �2�AdЮ���
�����i)b��eU<Q! mIh�u�%���CDh�ku�f̄Mr�i���su���T���3 ΀��1�R���<��W�0�Ț%,P[�ေ*V��O�=����zs ����/��mHv�"I2��s^۬V���ܑ�aY7�Y��ti�p8)7���q�����F!�aSɣ����@�y�C\Ƥ�'Y��&�x5�~��3h�s6��I��U8�8}d*Iv��"���y��_ݵ��>�{f헴q��1/��� Z��x�����Fa�dsڦ���W� �<����t�Y}��u����^�OxV�w������!� ^�sw"@�P�N�f�D���z�fa�U`����\�HrQ���KB{7l��WlK����S��ؠ�Ń�}\S���(V�'�^�_f^�g8}:��[�q���pSɓ덹�G9��҃겺�W�1e��K	��	��k���#2��_�M�;�)����5m�+\V�͘ߣ���IabS�d�'w�|��U){ጕꎼ��zՔ:�t�?0��<o@��N�SL����a�i��G�#!�8��Do
:���{ғz�gL8�)x��B�`D�C_�[Ű�n �\ۤ��Q�l5I�d���LZ$�H"&I���ֱ�=��9啖T�񩐳s((��X�)y���\A�W��a�7�[jk�N����j=?�Y�f�&��ۏGm��2�.����]`�ȧU�Q�E�8�,�]x{�켾�?��f�RK����?A�"�5��Sh�w�Y�0˃�]9�7��O�>Ca`�{���+�Oq�#��1�z��f�ki����]8�S��i��mF�c�����h�S+�|�w<�@v	�����^�B�=�P�
:e�����D���
��8o��ߓ2��=��u �W���+4^]�3��	�H�l(Ip���+9���?��8��(`����'���2������]$X[p%�G��_AH�����h�-�0�TN �jC0�7�����E���,.�<ԧP������B߯);!�>���d��J�5��rz�
]/��>��(�\l��#|�^���x����hbMEm����
�V*�*bjʗGw��R%�1��[��}e���q�V��.5��1
Zso�8�Ht��߹�g���oOP��%��~1O��(��&&�����9i\�$0ۺ��"U�ǿH
Ap(�ˁ-m��"7K�-�Tzwo����d>fR,n�fk�����n#RL�Si	T>�{Ĕ[� q��se�pY������!�?�g�v3�/�K�a���<j�H��Ey��.��w-����y��8�R*�aU�W$ �9a�p����&h��2z�t��?�����.�L�6 �7DN)+0J�d��9�8�\��D�zE�=�Ku�j9(ˌ��<1H,�Еᜏ�����I�N{����~W*�!��C� 3�>Y�h������cJ�\�A�B7�o:5C���آ;�e�d7�c6my�����χӛ���	�ׂnm��@�&�.Q�+ �C�^{�-/�啦����eң����f���9!����ˏGJo�,��R%��V>�2&f�>v�m '͚�ޫE�1���0�A�>��`��%>>0}��2�ʄ�k�"pHɄT+V}+
Ѡ�&�>�.�z���X���nf+F��j�#���%)M�l��U�ڼi�*�R%�(]:di�N��#S�NNݗX_���%5�����O�PݷВz|�M��n���\<c򧭷M���7RQ�����_c�7���_.$z)m~}���uc�+�0�ʱeC��f��b�l:]��l2��h𒖡�N2�Wy��H�YUg,v�95���]���Uz�'ŉ]��!qU�՘��L��W@�ga'xj�0��}|'p��W���/ݬ��AP�j���r(n�	(;�7��5��dȞ�[[���2n&��Uo�r�YX�ǜ̒x&]��D`ޗ�Y82���!Is �����A�j%~�1����=>��q� ��:j�j[F�{�+���3o8l����KF��,�O\�ac*�����8c�Q���s��B�]�5�h�dr9�q�{��+3��
�a���y��[�-�p�jn�Ы��&7�dZ�0��F/0f5�1-faɠ���.�� ���ÙⲒ]�_��A����x��a cWm���Iu%�uF��+���.g�d��[N0���qdbg��r�flkǋC�VI��{Y���+^�C�(�Ҋ�N�~a9y���8_@����&�}5��*�Sz(�f�]���Hߑ	c�'�z�C��B��>�D���u�/]8��l81��>��o!�s��B�](�f֒p�M���}�2���0{_�:e
��]:��L,]�4�۞|�J�'R�e���ꩫ"��pB�+�= =s�/��+�L)�![gC+�q׈�v��8g[!:x]���!��Y&���#ơJ��7��r��*mzx,�Qg��P�rd���_Mr��>Y3Tg ��`��f��5m�h>�e����hpR,�-�k��Ap�����D��'Ѯ=ǁγ�ϐ�/DC��{�����)9S�tD��>aP �G�f��(���]?mCǤ�V��I�i�:��*M��k����r��x���K?�/�Tl���B'��d��}x%���yRrK�Z<t���$_I���=u����B��Q̚q�bc��У�/��2+������Ei��]Y�� R�l�t9A�{Ą�G�Ǆ�%3TÌ0�=A�:�|2��L�-/��߇�4R��(`X�W��ܚ���k ���A�˹#Hqң0�8b�(X5��������\�C8 ;Ka(zh@� ����Uz{���!�@�Q2�;;�kq�M�5�E�C;a��X���~c�+�Υ���ނ�	�>��B�"&c���l��xY�)����}���&Ց��z\����R���@�"i�;׀�-���M��D>z�(�&����\�+���g�*g�����ԌoJ�	w��j�=?�H9���FmΎȼ��,ִ���M���V�>$�_�͊�5Z�
%A����gP
�V}�_\�Bc:v )��3?�poȆo�9����҆��9�Ď<��c��r�K��b| �� �>�<H����`�<<O�����*�|rz9���+K����C5��q=yR������oH�p�{�V�-�Hl��!�?[���56��0��P@u��rx&�D�(��j�|5s?�o�U�`�a뻔�o�K6�'?���m�a�x�щ9�Y�3��e����7#�����8������y�G�]�.�T��bG�'B!�2)L]/M���N�Q���S84���sN�~_��|��T\�I�.P��ԏ81�C��9�k_-7��HvZ�^����=��J۹Iq0�� �2�Is��N���+��!N^�g������p���ӡ�*O*3�5 �:�W.���ޮ����h�� ��冀�9�8vu���yQ�F�ɬ��m�n��:lB�Է����q���h�EA�B�j�K�d������;
��h��R�ѻ��,"R�Ӻ�אOwT�1I�é�V���\�M��3���R'sW���|xs��f�����~[?�'86F�����l����8.���S��e�Y��F�<Y� �+V�1p���HW��SJB(a��!/CZQ�RnjFT8���/Y�A�96���-�W�1(l��T}�|�v@/�(�⏗[V��j��<nD�Qquݣ���M o>yu&_D�&��G����0^��R��u�m�F�M���oL�FۡAumץu�9]�����ݩ�@b���b0��G��,[h&K�`��/|$��y.*@�yz�a�T���w��� �Fc�{�������%��Ӧ^�/韜UQ�|�h"}��;�+f`���s>�}-t���}sjYt���sh������w�W�Co_�4\�����,�ܚ�PT�S�Ɇ�+[8p��&6u5�Sm~�������R}��\m���D�P{0�/��C�B���"�z��\�v$_<�0�]A`�Y0�v��p���^�e��_{.Py��J��ᷤן�̹9�$�!x��ʴ��2�J��������w�yA/��-U?)fn����m� ��\�6�WS�h@V�@��O	���̘�ԑT%���W��k��0Qf�<Tՠ�1�f�jG�������k�~��:M������ �����r��pg�o7��NV�R���=��s�Q��*��=�JeC�a2�
��-YQ�:@Q��ò���U$Tw&�4|��j1b���&a��j)�z�.��hԶ�B��T(�O[��f�;! zΉXP���嗛��;T��N�� Y�w_���u��J�^Ě;��8�*3�2�
6�<#A�O�q�L���V��q	!�uƐ���:���"�*b}�
W������j�4�$C�<��n.���f��%��A.	�W��7�Ŷ�L��󈸀)Qu���a0�&jJ	�MS�����w���Fb����c���9=����|aΖ+Q$���j�8��ޕ�a��Z�f#f+,s���ns����y�剾V.I6F���Gq!$V"J�;" *14�.�k��P���T��6@���?�y��J5����om���(D�Q.3����K���7��E,�nJ��7�Vjz:�Ƃ#7�OSK�g��`�=��'�W�G��9���A�mT�����gO�l$�u3��ٹ�']'@T�7��q����V0WC�T2����OJ�ШsY���Y��G�U��ݭ/^���6� zɸ�?��f���!�d�4��|�%ʦ�BY��	12�ȗ�����u�/k�2�r��,���L���v�,{Z�D>��^��J����j�W�.���r�qc,ьv�{�^��ߊ�Uû�<�j*e�b= 6R�
o����2M��V 6���I�-'��W�4����h�w�e+�����񈑳��3�k��Y�;8����ĽE�P���X�
�ҡZk������	�X9Yi��K���f�Z�X)�G��qc��0��)9'�d�V����ԝAu��B/���<D��9*>~ӶJlK��b<3����V�V4x�$�j�4k-K*�oh,S�!O��"��*���r���㰆P��C���OD@P��3E�(��~Q��槼���;�i��KD�������Iz8ѓ�c%sD\�P�GQmq��p-/�T�{4�˶�T�&����H�Ji?'�λK����� "��\6��;k�4�[� �4��+�ەhh� ��41�|�h��κ�
]�ʟ�܊b�"�oq��|���`?�q��.�kA����n�ΰ����s�?�&*�#�o�?�9����zWr�3��K©3JW/���Q�����������^���ǹ�I4^	�]��jTY�f�y7:hk/��֕�	$�^N��q�c~Kݮ.��4�mCh{w��<�ߞ>4,��i��*͢L:�p��CII��{��V�Dp=�T�i��.�+���mUc�ߞ�<����ۀ��E�6�AL[]���Ȩ��5	Q wj�������$Ԯ{�G��Z��x��R*	��$���uBBNa��ǆ�~�Kum;�k��ڴ^IQL�מ�t/��o�'�E�Xp��w\ł�m���M>����� �)a9ۆ��0�"	'i����Tu�s\��%O�Ѣ%��҅������5�9��4�ՓWl&��������Ov� g��9��Pk�P����y��9�V�_m���":��g#`g�<���J��oC/���JY�7ڨ�9����㈬��7��Z3�i[�u��������5n�>[�o�p��W��1�{c���x����Pq�²y�\��"�4,g���0�)�I"����z�n�b�I%�pd��{��K��Y�(k6n(S���05]v،*>r8�^�����z��l��
 ��@8��c޸�S���>���
y����	�m=�l�MZ���, �s���'�p?�w���Z %�Ԅ�\�U��lX�|�� ��"r�~�Q�֢�t h1���-�]m@y���Z���������Y/�Q$����.�=-��(��X	�)�q�G��dm�V�6+H-[4j���2��:.�V�0�.��2G�E[D��I�zp#�%���
����Y����7<X�M��5A�y����$u�&���H�&�k���a�N4#�g�	8�����k���W_��G�`�:z�F_�"����vnΨ�Pc�h0g%k���Üy��(
n�3�R�;e���_�acw9l����p��
63�u&宏a�K'758Ɍ��U�+*������D2�� A����@ݚQ���K�@��e�{��1m�\@ܦ����������)f$]7kw(v+\*��<g[߼S��*��w�\�����M��������o�I���S�;��7��8����^�<V�Ѷ׊���R�g6G4|n�GDl��լ�y�k�Yz�`��ӆw�#��6��6?���������7t���"���e}
N�hɥiO}Ӳ��V3��o��wX+��H}.���I?k#cfg��d==5�y���6�y�����Ι}�MY�d߂��^{JziO��5&X7�N�-��+og�&}���,ۦR�Η�6Lό4��پ�8)9�`l#���=����j6D����p�T g�.�q�wy�<o`�tp5��NbW��O�-,��gO�����\cǛ��|2:7a��TӚ@R�=�����$��Ķ�HZ��!s�^�~A�s0Y���0�#<�h��ڿ�j�����nK��+�s�2�抙L=7T�A>̛��f5����8��k'��QkU-�4��
�g�O���������&a"�����l7td�:2R��Y&�2�^�janL�0f����a;[ܿ����&j����7�w8�ÔFS�5��+|ĄC����M o��}��7��F[���|<cֻS6"�L�4F.��w|����>��-�:��0i�����d��Yt��u�1��Q1���/�^�a��u�Ψ����wިΕ�/��};фX�WJ����ss��l��7�;���"7m�����*Ϻ�ʺZ��b�!Z����L�H&
��<00�k����Ġn�)����d$�ڙ7����&E.�Bw��g�Z���>,$$/�Z���>n{cF�DJo�Չgɵ���W��e�M<[u�s�zh��T��N�OdT��d[�C���R(?*��5��?����F�Q�1�M&��W�_�!��ہ�-=�}*6����w뺅��B0�J�.���vd�����n��n��"��	�̗/tq0;�+��L�*����Mx5TA	y�\���~_#�,~��"�/e��4� [1�����=��?�'(���4jV��~������'�tIt��P�c��^�C�V����6���S/ �a����m��ZƱ��KM�DYr�3�=�����-;�qMK�7���#TR�,Ml�71�@�LV@k1F���Y��m�g�<0�^��,����$��HCW�馮QtXQ��e-	�& �Ԩ�tSk���=!5ö^eT����Yal3��ft)9J��
h�ޮɥ7�.2ɴ��g�2���㠳�Bj��"��� �,{��/Bu*���(�� n�OYJ�;�MDlx���/3��s���E�ۡ\V�ͦb��|tL�t������`|t� g��6��m3���L�*��V����.7D;����mi�\���VfM4�Es�!S�,�xZac{����t� �ɰ�6Q��
�����AB��?,�$������t�����X���,��"ۖ�`$]��Ál�F>������}w��f-|�Ep�\�,<�8�U����N��5^��E91h��=H_�Ud���i�bh�7_���e���<�B��M��ַv����6zH^�ŐT���4c�jt4�x���o~MG?��?��9���@vi}�Z3Te��bJ��v7����<2�2�6�2��)�/�B���ED��t��U%;�;�j}����vW �Gbm�4E�2��N��b8��+��G}��
L9�T�|KI���m6��Ћ+��p�^1pr
�}��`�!�a����a��Q��ց:d��fGac�_td�FbA3_^�x�(�s�����T9�:� �5��Ass*Tw�+�o��(�����:�6.vi�P�%T�vuD�(F}�k7�س<�n�-1�̱��:����$�]r��:xhHa�a�@�X��N�vKW�y�|�Jڨ֋F@|�>B�ɱ,=lf�V��Z+�!O2�����g/0-�/�/mZƏ1@����x�FZ�[��>�k}s�T ��*��«���2�S�>�G�L":�S��]V_�85�{*�G_ǯm��f�	?�!H�����cQ�'a��=Ѥ��k��S�%;;�z_�&��^q�/n���;�kz~HSA?�#e���s���*3uRq2�D׈y=��,U'9�4T&��-�vLmظ�>�IԞ�̀�5<&"�=%|L����8�`�w2;�+� �H���pӑ�NЖG��(�N0$����� ��.}�(cd��X���I��S@[�h�]��v�풲�ȗG�G;�-����Y?1���9�_n�h��C�O���7v�����}%�^�f���E����~L2�������'%J.���E�L�X����	8V2G���s���2�SJ����T�F,��|3��=~!�(��7hEf�0�;� ���P��6"+F�GU|e��@�u��C%$��b;��T�<M �5�_.|h��HE���L��"ByO+���)������l��}4�n����f]|X�p�.�?��iEVHG7�KW�w��5� �����.��P����m�����7z�dU�u�ڈ��'L��>��Lx�+:����*�d7�]��6�gySl�ct+�����U���X�;�OWW�hG[��
�kﰿ>6��[[ob��B�h�K���P�w.�M�\�q{��ID�,OK�bB��FI�N�x+ı��L2KRd=J�:�m%Q�;Р0$�`��&����L�z���@��F�TJM�Q��2�[~�$�&Z�#[��wZ�N���}��<�	��׽4^Yhŝ�bI�ƪ��ܵ��; �d��r'$�T�7nᗸ	����,�;i���޶��w��v�Ȫ��j���[��wHɳi/#�B*/��'����E�JU�2yf6�W���[3Λi�=.
��EH5�'������;[醮�EV��
��p2x�(
8� ���[����EO��84��R�=��i�wb�	�<s��Z�*x��r,ͭ��ZQOO���ٹ4�nnhJ>�+�`<-�fSjnP�;��C� �S� <y�c�]j�(��6GQ�W8��x&gK4�b5���L����Id��I�:eF_/[��M]��������V����g�8��)0*�����#����ۄ��߬�#U;�.sU�O�PhO���[�� U��p�O9�꩒ҭ(�܋�4V:ط�"F��Ip"�l�e�$�:��3��\�ϨV[rb]���<3��_ ͽ77WQ��#nn�:�>�аk��@��ڲ�5՘��>paL,x/S��	@m���d��?4��2Sg���*&~��xS@qEʝ�>߿$Ľ�?ɷ���.L�5�B9�sun���m ����|Ƚ^�FsjCP�-��Z��s�`�*��w��@U;Z�2�2,�f--��<���<���7^�+���y��{-M�m�iA���ܵ*�`<g�2��t�X��k�Q�JF|*5y�A������V+{�� 4�mH+j�>�|���%���m��V{���$h�O�<�@�Sh���/w}�(��T6Z�t�-E�ͷ��|���'�&	�� �	p�&j4�y��`W�u_F4���V���ab��b�����Oa����:�|���T�,9h$�����ζb�< թ@����>��,��k�M����ąոMiv	�t�ʵ���rQe�|z��ZF�?d�/y�/�6�/<҆��[�k�7��&0��)wc���	&�Ɲ��ڂ7������<{�&Q�������.����v��%���iLX����ne�3�g���OF<
���̈́y-�L&��S?c�/(��p����yMp��dc�J����8�Q�1�vm�O}�y�$%�R�ui`��ym�W7Q)���ke��(7�:�����Y��Nsq�+���G�[h��9�6�[��|:���;@Yz(�tu����f��%<"��ј��e ���5/�Ch0�D͏X���V�Q�������s9ly{6�(���(����D�n�.wQv�rU4��Hֳ���hƹ�|��/�?Z~�a��=H>'�]�tL�!@��P�T�W�'�[伶&u^G�PZG�J.8�^x@7�<@�~L~�����)vd���db�.6PC��p�����5�Gȸ������.�M�H۳��P p������r���I�z�d��!�N�.��~Q�!g�+%٦���z�^.�� MY��o$�#�d�/)��)��
 gj���^,|?E���3-���ק&��[&U��-|�ϧ�Ç@9���o����n<�ѵ����9�S��/��7�1D��I����(��'����^����Z��%��"����.��K���-\h_6w�OA1�����7���Q��6��F?�Y��%� Tih]�v?=<�e�9y*(��f��,�Ơ�?�V%��o�Z�� Ҭ5��|� �����'j#��(�i`�2��s;�?A���� |5:���������.1^����x�_�� �om=�mj4����.�0�J��E�}�����ϑ�^K��h&�{)����*���}B�q
�E��c���Ğ����᪉�M� _�*lRy��)?���,�C��e!=!ȉ�9s���H�[q�U�1���)�9ܾ�?.Ǆ�"�Պ��-§2 '���f���*va�8���c�@�,6�
6����ׅ�s&[Ļ��4 ���qI�K�߀\��B���<��c4�[��9��r��c�x��`����V�w\ݫ�0;7�s�R>N��<�c#�Mz�
#��9�(!-�� �Kd;�X��ʫ�ݏ�cWo/}�l{��⮿��Z��!
��ְ�J�͸I�����E}��SD��%�ݘ+�Rn�P�%m����7ۘ�3p�6�?YT��O�Ɍ��HO+��9������^/�Tp����Am��>�����Y���;�C�$bܤ�wsu�F�D��Ԕ۠�Z�,�Y���EF+?��|�b�p�
��3���/�ᡧ���qB[�Բ��S��I�R��b��4�xp%�᠒F ��_
fJ�qXut��~^�yC^z��X�E&oi�r�z���[d�M���`�{j �EIf�>�H���C���A,��e�?S˫��וmZ��ѱZn�/wr6?*?8�g�����N��������{���6�i�2�Wd�G��V�jع��c�[Da��ة�4L�x!0
�Z�z{��v��W�=>p�Qq:y�<�*���s�/�5CJ��=���YG5{� *e�0���mR�qC"r�^a��&��[@≋Ṉ�,�Tw��:yGԯ���\j����Ώ��~�?�q ��|l�WVB���|=�X*\�yǺ��ŉ5dT|m�-v�M���V�n��{p k���"Ow1E-�@�}K�Tѫ�L`x��f��$"�c8��g����Vh][ӜAJr'D*�rq���e��sB�w�:Rgl��Oל���ƾ+>TWk�����QQPh�*G=囿Czcn�6���x��+��s�&��� �U�"�i�>Ѳ�#�S=ōG��I�|O%F��<�p�>w^��su����s@�°�������$~+@��Ր���ŬP�FM�`�=Nf<$��sD�?[l��jbǰÖ�)�D.��n�Z������-	ig�SN0�^S"ʯv�ht=5sD����5�H
���|�_e����S�@���\��-cIǬ�ɛ�Hӌ�I�3�O;>����9���X�7X������ꍒ��!�I]�#r�Lג��M�V\�]R�QA4��s��m���!y���M��O�۴��a�����ƶ�*e݄Y��GB��:4'���(Q���jFH1�^���3F���&��/�����K�$��-��Vb\	ߒ��@s�ӡ��^��,4��Q/�'���f8�	8�Z!U��¶��̼b&7�:"E�k�v֖���"�&H	+����3�`���Mv�N�$f�0��Me���,z�&3&I^c�R��К��C[��=��/=c��I\���(J�-�Y_J��Y�(`e�N�����0���];� ��������0���]�/[�N	�_QD�-]�i��A��Y��$���Ҹ698����Fv�ߣܤF��pm(�yM�����xLq�G����m�*m"��$��=k�AMv�>�?T'�O2�	�,�K��ũ9�D�ױ{3��CW�L��K�~���=U�-�/�Z��g#H��ˇ�������\;P�Q�zՑ��Tc�^��q��7X`M>]�8M��� H\e���D��~�B�-�U��$�_����3�d��U]��l��_��#(�����~+߆b��F/d��$#֒�1-���֋@�ˡs���F�N��_^��7���d�t�|�w�S���I� �R��~T_ʾ��Ik��O�}6���A�G�o��ӳ�_�Znb�@��2��_Nԑ	���^��P���Q�~C��{)�QX����s�o��ezy��=54���t��>Bc����K�f�&�����h3f��?r��s�n �m���\��v���4����Ə%կ:\�}K���x�($�L���'�n���#�^�wi��-�,�,�a�7Ș��Gz�f8<_�i��i�/jZ�Jm$�m73g�=�v%3�px�ء����/���H�ԯ1SvqbM�/i`w��n��w}�<�f"d�����ȹ��g[��es�Lez�1}HKRE�ǘ9�+7� �'w� H��6c�j77����!�l�Ո40��[{\L=�!��k�7�Y�˦?�l+Q���x�Wi
*�i&�^�j�p�v��4K#���G�[%�p`�ą���깁Z4˿���[b�&�����������<�`02��v��H���	�~�G��Tp����c���	�t�A>�f8;��m��UY5��?XWB��u ��������}2�����qB^� ���2c�}VQ��m]l�9��v��N�_�=���.�PȰgy	r�eB����JKnHG�%!�Y��
n�����[���n��q��1�nM� w9E�BS�k:~����* `|~|���=��f����)"Wjɻ�����9p���0�`A;���(И��@V�G��h��!�����2>1S( ��lj89^�/Ͼ�ݿ��.�V���+�����V|� �Y�&�����!��H��v�6`20D�/(j X����Z&xMr�?��*gf�T!4���έۥ�-ƺt������U���55�Y��ʓV�A��t�<9_�J��1Ed�����\
���D����n/��JGV!��� ~�'��V��>���k ' �~s���s�O>��$&a�w�ʴ�����`�g"@A�m'�2�Uq�Y�>���E���
���P��g�����#����J�u~�Nt�����W�'�&�(��|�|g�w�"O�.n�k�ؔ�y4�`����73��!�C�Q-5$�p�GW��(��[-�,&�5��z2Qt@>��B���T&��!��Ή/���rLz�D�T�{���d��?�O'�� }�cî��9�hPj�c�s�ӝ�Q��w'�2�@�#0�w"��#���[d�%��*!��"��2�>Q��Igd0I�@O34�cPkJ,a�&�g���Vq:�oM�ʀ���.'�*�r���_I[�r��&�B9k��}�ȁJ�6�SM����uQ_�2_L�{^�(p��*�����Ήm�J��jF_ql��g�Z,m1�@"��!�T��e��1mH�<Hx�(k��E�k�,��_���A��#{��ɪ�Ἰ����;c�Gr��[3q�1̷aSn�~���'拖V��+9�A<�8��v�X4z[ �I�}��\�2�Z���{� Y������Q�^�ұ�4�e=pr�d��]�X��)r����l#Nl����)�VU6�	мu���m��tվ������b	���U���m~��{����ff4 -g�`�i���m��ǥؙ��|�Q���Y7(Z���eӵc�������Pg+!���4�ג�؏31�(~ܙ&57�a}�B����̢ � ���c�k��	,�E�C�*��`�7�7m���F��傞�>V���4��h����
�?6�
���ڑ�"�m����ͺ�H"����2�s��F|�?�qwuac�^�M�|/����4�،D�8⤝b��^�Ϸ�^��6��B�-�P�ckֽ{�
����������Ch<���q=m1_"���k˧p��h��=��E��~�As-�:~lz��6}C:��t��+a�f���:����!�,�f��K��6nܥclEp}��Qz�̱g�������q��W�,�%�".����Hrޒ�</�TW�O��ޚ�3�=�����-����<���X�& �
�׀�τ$r�!S�v��E��Yl�=���N7�c��$������(�
I:�K'I?	��V����2w�`!kp0���r����r�͉{���uMs#j���tH��Xjo��r��i�!���ՠ�iq�����ܘ��gz��Vd�4�xK�,�B?�H��<��	�P����j�J�U2,�4_�˳�,�"���_�ӬDCōS-V�V ���n�ˊ�u���E�f3��b��j֍4��Z�ہ]�Ңm��>0���Ofa���Ȧ����͌
-�T�*ޥ��N%홒��L�e�j�z�7�0a32�F���, ǟ�j�E�B>~I~;�G��L5�2���Jޟ�TL�0����fLG� �}���1��=āW�-$d��
B�d��s�-E���-��#��pyp��H�]��V���R�n7E�Ob��XQ��P�0:���3��ƍ1㣂&�v�g2�F�-ӭ��s�Ir�c�IR�Y�z#�n���C�F�M�tR�K�� ���� �P�n@��i��q��;�� �@.�~��q�cW�XqtA����@�:���<l��ЇK.I�R����_�T&��q�s'v��h����P�s
	U8�
�:�nP�%Y=���Dr��oOZ�br?��D���nSܗ���ʘ��dx5��Ph|�3݆��d:���X�׈��6׎s�4�C/��;��v�\�E�!)�Y��@W_�l����w~��u�v�,��8�UGm&6�N:s�"<��k]����gI�h���Gt>��F���n��M��-�X�z�b�4���|tc�9;�4>��%s�>;0������J�gr_��j���m�9u��q�f�����1��A���L�n)58|�d#5���HAς��"A %������Y2����,I~�_��t׷����D�l�-�XģR�d���-�`�2�I�B$tH�b�3������&�=��Ts���,��pb�I���xOV�
��q�c>�k�b�\{ٿ�?�ubHN/Z���b��Y�=޽��Hg����������{��T��v���p�th�t]O�6D���� R�d�^5a�G�m}�����!�R�Õ���/-�H��['�ѷjJ�Xf��1�!�oL�}��E��r����W�ll���a6�ѽ[��B�������k'�¡�߳Y�`���Q�\-6��M63�Q���J��y��c _�ЅbD��ڤ@H+&Z5%�����w�>pAM���f'��,d9<�fQIt����Tn�DnJy��"h$#�;~l����d�U��!���my�Қ� YDgK����g�6 [%H�֘5�����ˢ�iX��d��#��N�f7j�8�9!u!`Ў��@~��x_0!�����cm��_�L��,1�9�gO,��*�+�R���U	
������8�`Y]U����ż����A��,���Os��B�>e��#��43�n;)w��������{��$u�v��4س�'�P0����ڵ�.�\dg(��<��ANK=��J�"�FJ�h� mY�Y<&HD#a�gW�A���_�>�/��[��I��v�<J9��r'��Gr[Du�5��M}̜��T�OK�W���P�B�P�2���7��?��|{n�#�bG^(��l�?2��(O��H#�P\cЇ7%
�j��^�u�D�w?f�K㻖H��&��:��pҔ��2��9��8��p������3c�C�Pw6l�tY3O����f��)�<��C9``q9��@�f���)KD.3��h\fm�����dT9���fǞM5"�d�ɵ��=Yu�F2��L+�AkFp�`c�X9�L��	C#�u���@u�Y*�J�o�Yl衈��������
�F|�EӣD$B;�%�ͼ�ϠOz
<)�j�\P���hI�X��|�JH�/ќ�N�xD��8-;��R��J�P�f>�{�BN��
_���=�ƣ�;��?����c���RB�M�N�R�O�.$�������߬p���30%�*`�4���|c�!9\���c=n�L��H"�Wx��I�� ��R�=�b�os�/"8�m�!�X?��twu��ӇS��;���'A���z6�	t��2��Fw�=S.S_�g��12���}���ɋ4+'f�l�p�wA��8X��x'b��l�({�7�z\X��$i�43-4FT�H�R�)��sǙ��6J��2�ԓ�`�H�P�6��R
gC󠺏���a�K�D�-��,pa��ϡ����<�Mm�TJh�9IQ��f�N�ƿ���g~���i�=���b/�{�}�"�qd���f�+g�Qq_�P��k�gn�oJ�T8������A��#�D̴��JbW�%��B��(��Bs��R���g� �5����:��}[�VwӿD_����j�'��V��5��&V�/},$*HS�NY��	~��"�r�'q��\@j�]:M�eȰ�"{�5:5���VCM")bc��'bs~t��r������E��e嘆_�9��-*N&\�ZN�+-�5Q#`^	vg����Ȁ�n�r����q��-L��g���y�94f#|��Oz�Z�m�����+"A�glu�X<Nn�˂�]?���v.x�ĳ;d�͠���a1����e�	|�Z����ԭ��t{��Ɣ� �����KL��G��I�/+)��gH������~�ZG�ܻ�+�3wq2M��h�ĳ�����҆E���Г�>o��e��kp?�k6�F�4���D��m�
L�q�y�;�o�fL�َ��<��j�u)P7.��H|��Z��͸G@��?b.9-uM�������gi�IM��-���G�y5������#����!ڠ-�7�}|����ghY�1=kƏ�0\��C����

���;���������v������EUÆ�����2==����Y��6%#��2M8f�4j�!�8@��n��Z[rz�P������� Ŵ�%�N��{��y���,@z��:�F�I�'R9�=���I~Fq��6�1�To?',�|F��v{i�݇��D(�$
�nҠpk`��k�޶����������o����٧d���a0�`ͺ�~F�K��@���^�oU�5}@�#a^���
f���x�?|X���s�Ji�O��� �E�9u���8z�U>V$5C74�Q��������X~��u�8}��rw4K��W���mnXֶ�m�������L`�ՙ��s��g@��Nr�H��X	ii`��3�۠?@���cd���=_jO�m�"pJ8Bq:~�}���"�jhbSo���:���)�[}�~� �$�nK��|��#�˕�I�����M.N�zN�6��_��}E/tPy�b��oð+��D4gS�S�&���.�J!�5?�\�_t'~S�q�7w,��s2(9�<2 ������B%��c���Bp��uJ�������%�C��?�W&#x�f���1̳�Ya�|����^bִO5g.�چ7X�!�Y��I!:�f;���*�W�ܙ��W� ]5P����ܘ}pg_�:�\f>^��g�N	�X�ښ�~ZR)�=T'Rm1��!D�N�909���.���ֺ�/�;4vǽ��ܚ�ݞ^X�W?�\�
�V�S3T��������d�h�
}�
No-�����p�~���nG��0H�d����s�
���N���ܴf%� ��C���:��P�]D�r��6���/�+�ޅ# �5II�[��]T*J��	�='hK/t��p�$81����\��W���c���	¶=��8U�hg��{�R���_g�1�n( H�� }ND���eϱS�0_�Z	�OP&]#�L���6c���w?R������?�`�-c��Q�����h|<��j�L8�,2d£+�p���`|'�:���U	[6���V6a�`d�����J&?�d;��� q�V�f�욑Mr�	Y�d����q�c.����̌)@�V8/WX�����cU�V�8�>͠�;�id��|yͷ�'6�q�͛�@�)lju�����Ԁ��14Ki�N`��P�"�PZ�Q;j(�;�S[AP��ŷm���rs���n�΍����s��&�׵?��\=t���)?�	��V��R� ���D>��q��'k���ݭ�k꽶��W�����e3���Vx���}�M���P���=E`��o����v7�{ok���"�KTʤ�5�X}����Z�������U�2\O&Sރ�?Uc&(��p#)�k�P�Ԕ�����,5�K�7#�m�6�w�AL��'0w�Cs*�@"2���4�p��^�I�P��ԙ1�ī��;0!��������;�?E�W��ID��cn��	�g`��Cڶ�)C7Le݃2�����4"ĵ(r�v{5�:�1;e�>���ssګ�{����}��o�����Fʮ�řK<Y��z<\�T���6s�n��#+������/��2ҍңd��JrD���Bc�!�3Q�����I���Q�I�L�|�qw��f3��@g�`�u:v��]A����.[����Ѷ��E"��Xm@U8`��Y4ꡔm=���T�4ht��SX�bu�B_�M���z2+����O�;��×@F�����	�}U�
����߇7
0S7�B�}�螴g��N�#����E���hT�LS1�tN��7y#�[�����2f��b���B�_�#ʶ�2���;��"�V7+>��l� LEFq>�p��C{���2S��t�uK/��硳\���m�����"�Kj�Fxt���Z	ȋ�b2������\F�K"� �3as��Szc��@��)d1"
���2�R�ĳvZ�9�K�녎���п���4Y��`Pc���q����ST8ٺ��O�T�Q1@��m���Ns4����t�}�I��7�`��Ѣ�V_�[X(CP�����3����&~�P��Q���$�2��^��|6(-���-5�ٰ��Un.�vĴ������"u��~ู"���a �_9�$ygOY����*;�"�95x��4tƿJtC�J��BK
��������� 4�c榱&<����r1�=�� 6bٶ�b�t��dK��XҠ^�s�*8�ϬUDcGbE�e�*׋��(�����rϜ=C�ћ�Q���&*5����u|�y�"�vwJ��z[Ɋ�mH�t��f�3C5e/~D~Ў%-�
�|&z6%��Y�ܓ�A��w�z~�~�}�:�H�ӡ��.ȧ9�SZ�zUIn��os��Q?"����a��/T�7�o�q
�F�:��ߴ,P/��������a�$��R�΅`��\8���)����)�H��yn`(��*?�Na���-��f�F�W�B�f�Z��ap���2�4v�_`@�H�`.n*��-V���R)��M�	2t��з����^k�W�Y�Fġ|���K�$c��x��@Ln= Lq,''�`�0�j�b-�#�P۰$�X5G�Ez��4!~ƛ�-�;xS��� .r'	_����)T��lݠ���1}��.�4��Pq�x�*O�W�k��!i�/=��^ld~�����TzS۔C־��X
��(�eO6R>K���qT�ʩe�$L|�1TM��sP�7)_�F�.�BA tt��F��_�Hq��!X�Hۻ���6�ǯ͓�2�ǌ�&K�J��2PKd����$��'�9P�+� ����>���E���$���n�*$��hT��?ğ��ŏ���T�d�_�.�6!]	�i�6�yj�z�`�����_�J�K2���	��G�DS�"����2�K�+Ff��l#�����ܪ/Ru-ƨ}ݴ�YBH*ٕ�q_=#��g�n<�N�w|>8zvX����F�\��9(���6�F�m Y~�����3�(:����omƟj򟎆��ۆ|+�sa0����Pt�3X�Q�����SR�X������/yL����8��8ַ#v�#�%�r:QY"�E���1]�Ӊx �i�0x�tύ�]W�U|�v�Z��m�<{��7Չ@���h|��y�`�0��,�DƠ�*�aՕ�N]��L�!�f�#�	,\Ϻ>��g[�����e�;�$^��ժӆ��>yI��
�:Kk���Ȕ���)���#�s����A8�Vh��Y��A�:f�@I3�*���-�fh�wR�QgA���r�C�8�h�h0-5��3�]���]د�VQ�Mhˣ&�o����7�!u4�j��K�w�/�x$>h�\I�#�"�՛n�
ZۋǾW�!;� �;�*�j��&�;&ډM�@�O����)�� �����9�I�xLJ�!
Y�.�(C���nyB�^��U�"���u=���U�<_�f��|RL���a�jeT���"&���[$�:E���9��ɠ�z,�#��#���J���iQ_�؎�V}�]�^��mO�O }��#�qR�ks�����'�B�6�ʌ��ɳ��L���~X��,v���V�j�&�z�-�����ٝuR%�����9������K�/�����u���d��*˺������#W�·�p)#p��͂���H�0�r˪럳��4�Ms�� ������	�7��-s�`�{,1���ΰ�1�g���E������k��)�e�����fV��]T7ۊ�d�᧟6�3n�.�`���yN����}�WV�mCj.�����x�(�v������Qh2���|"˻� ��LBvbؑ�˦�m��2�P�.��_ٟl������83h���$+��-�/�`��s����"��p��y��Ʋr�Y���v��qy��JU�*"���]��w9n)���ga]�{{)
��|�&7��?�;�I�]��Gx����F�nL��i󇮧\��2Ă�10�ӵ�Rs�f0�၍��`���H��$�SM}:J� �����#p��~�zh9��UpT/u�N��?*��SR�Ma����m�y>�hNݝ�'���M�y2����}�JJz� �/ c�O�L,,EZ��?ߵsQ¦��� &��(�zSH}���w��x`����c���\,�h��Mʾ㶂Of����;��@�b�?/���T;�~8N��GBT�G�`���&�1ƏƼ���c$喌�J`�1U��}e���e��,՟N�����f>"�{�[ƅ��D�/*�-���Pfi=ɋ�j������K�um&��\��0)\`��`@��~�h�m,])0o>�Z��h�5N�����*C�:1�	��k�7zP�?�&�J��>���T��V��"R�ۉ��,��R$�N3ɖ1B��Y���X�q`�6���W���G���Y�U�_z���,��7f�>����Z�x/q�����f�y<�"���K�E�<)M�_y&/�i*D__��s���1K�'b�D���C�E�פc� bVH��I�<���r�d�[��`��)��:-�=g��(<>\�'b���q,-�X�@�TVg �^qkK�"����ԙ�_Qdཿ�b����-���.��@���+EAW�9kYE�#6K�Y5��k8�1�uZ΄R����X�G�v�TNY�`ą��qKrɛ%5b#f��ׇ��0���r�:� �LQ0_5���=s�i�����$���P$-I���x0= UL_�/�bEi�7��yo�z���\���<�ÚiJ��F�昏���
R��D�B�W�t��)���ۄ��iگ�c���`��;��C4�\l+��Ҹ�F�<�@RR*)u=W� t�T����e)����6q�Xv"Γ���E�w�~6G�%;4oV-�]\Z_A�}d؏٠"�4�V.�G7��B��t�Qɕ	נ<)w������#���R#*;M��bZ9�)�@O��·$N�I����Og�u����*�	�2�[��)0�w��[<�V�H�h=�T���I�8��zڱ2��s+t}��I̋��6���3΍}/�q��Fk{l��;ŵ�SEU*�N��ʕq5��!��4
5ZR����cY��|$h�dH�q|�A�	V��j�R��eV�P�pɉ���[l}��\��1;ޅg����;����l9��v�F�3?4/Z��y�>��ߍ���k��k��3
C9���q��!`�p�sD��J�쫏�K�a���.6[�aB��\�m"3��d�\r��������='���v��!�<jVq�o����V�Ա�m�[���Z\뷩�/��[��CwȂ�:r�.򯳹,�5�'h�lc#����$Yf���*�Ǩ�!5���ƴ�tdD�4�0d��p�֓s���9���]�*zL�������Ȉ. 2A��GY�g���'e�\�<x�0���ba�2�u*�*Q�n�3�K��D��p��JgySQP�H��v
�?3�S��3�F����~d͚�l�̷!��G����i�G:���Z� 2���2J&��m$
~��C�(��Ē�8(�ٷ5������h���)y�"��c��"}���HO�����wC����*֌xP�9�TUK$Ft���w��Nw[5�"q�����}l�1H�(��R�k�%�����%[0p�x���`1\m�6,JV: 4�p�.�)ٻU�z>IOkVi}.����Fѓ;vJ� ��J}�>
�Xٚ�b�k|ԇ�+~����^��|��x|�Ǵ5�Vq����0��G��B_��R98���[��Z!�ƳN����H�7����Z�R����ʷ��I�8i�b"5B��q�g\��}���)?���ޗ����ͼD]o�	z�Pu�ڑh���:F�"��d5I�J�kmő�e����4��[��fU㵉�y���j�h�5�rdV��engCئh;�{�>|����{v��iH�N���w���a�
5��-��k�f��~��u���6*�
ëS4��S"}�����W_��P�zXk�kI�KKg�SD��A,<�4% טA��,��0�C5I�����[���>�Lݥ��:%�� �r�}}��+G�?���~O�<jtn���,���]�눫lR��FK�Hm9�W�H;�����B��ma�kR���*,��Y_�	� ���Ry!��;�$�|����f��)do3��]g�����ySQ��&)��?6���������~��2X�b�8���uS����r�~_��|C�f�w���z�A�t@�:n!�%O��V��u]J��������U&��5�-�G��M1���9�2_�-��fk���Q�38as���mK_��F諢�XU����e�l��_�G�_p�>�I�"@����o��mP2��\�K�QJ�k�&��$�����dX	)9���@oq��7���t������a�`5<nc� �\,o�Xe0��Y�uI	VU�����-�Tځ(JK�-ax����(�i�}Z+��vgf�5�3L��#h�<?�`���tk9J��;w�u���K~i�O߸e��"e��)�#��V�"�kD�NYƯ+,vj{s>;���F$���:��&� =��j�ܑ��@~�&�Z
L����1��hP4���pT��fk������$?�}o��T���uuLx����1���ü�>v�ץ��υ�R8伩k�v/�g��Q���L~�4i�"��UL,��N�ZR`S}��#�6O˓���3#cY�� �3#[3�)1�Lmg��Z31����:����	^���%���9h:~҅����������)脰����&�mNP�le��<�ٽ�E�r5�>9�Ht+Ν%��p8�lVct�yҶ�=��;C�J��Y��-�:�f�/�h����}�ÓW�	`!v0�ǝ*��,u��մc�Ԙ��)�m@ż�3c,:$���L��,r�!��[b����):��z�����Z��L$��r���4����5Ǒ�?���L?�Ĝ�N�i$�X���^pJ)���j������X�:"+�}�4��?/_�j���/���f8�aJ3��r��:��4�)�����[	���@�Ǥ��mgQ�%���Z+�6�Lx��3@z����p�`R�.�1)���a��|oɟC+����;���s__�rN ����Y��il�+[�"��h[b0�|-�L��Y���p�+l
���E�*"�D0qj-2Πt�x?[Tq����Fja7<���yI��G:;開�h�|SC����v�j��O�`V���]�!V���H�b�� s�55��0�H�8�~<:O�pk�b�i���,Y�C�w1�+�g�
F0�0���}C�h�2�C��j����IK]���跚4����<��B2�1+ʵޢ���^����;"P��y	���`���3T<�4��0q�P���C򒃄��7���'Aaxpb&h�J�U��f��]R���\�L!3���� vw6�����ת}M���B�� �,��L[.P9ѩo��]����R��+�	��&��r@�کS������Q��7L��@�
���ɼ��xޣ�z+�fC��OH�<���4����-3��������s���T
 '�YX�U�C�Og$�{鴙� � ~��
7���d�0_C)�/įn:���8.���a�9B!j'�S?��x~��h �������DϝiR�V�&��C�O��T8���N��m)~��(d���j��k2�^��9@[��Ð�*�N���v��}H��[��-ƧU�ȥ2h����J����61B��U�P�w�16�"�$퐝=k�t�C*��	q��������?���R')5µ�R�H���q�rq�j��v� ��s����f�vfȗ��OV{#�Չ���k�������ǋ�s�'�]@� ]Ô%�cLAU��ܪz��_(Љ��{p6��#�(`�`	��L�0-'�=�5�nkK[K�G��|�l�vjejz�|ι��^��!�u�ly�6��L�#���<��a�YD��,Jd�`'_u�>�W�V���w��*w���7��b�1�n��_�h�`��i�0��1Z�c���Њ�J�@�x0�[��F����X�>G�^�8D,®8��*�N��=��iHX쫠��`��u ��%A�ʣ��i�O���ϒ�w���Ȟ��
���Z�[:�Kx�W�BE����f֋�^�	k��)��(w������X��=q�J�80���<67��ڡjC��ԫ��f·ԧ�w��8������&p�{���[�!�ۓ��E�$���3��ҷ~���Y<ݸd3+��8�y ����O+�*�u(e-'�s��H��ҞK��+J9���|}��M���tE�d�����6�Q���X�d>�Ώ��IC�Y�!E����Z��~p?�/Qw�j�Ha:+������Ҕ$��UK��7RLJgX`�cL�+J6���~�$8��F��������vP>�P���r*,��(�j���/H�>^P=�h��g�(j�{8�$�������������*{�7:�0�����bx[淚U����s�?�5p�]߯*k&�&�� z�W੼�����s2����N�;q�E�ML��6ۼ)A)Ĵ ���6�A{]]��Ă���%#?.��/
,c��,و�"#�(g�t<-�J���٩�����\2��g�>}Dg�A������R>};s����5s�y��zy�a�^aP�����H	��O��E2�}��БAZ��D4h���p$�7����ƻ���ҩ"I��]-
~<����\/l��Ƿ���]d�=��I�l�TJ�z��}!��'N�JZ�?��������w҄}9@x��H���Y8� ׅO��lXv{���|RA���:�ݾ�@��)�is������
��M�:�A��p� �ilq��M�*$L�w͹"��SH�d~���
����h�#B��S6�G�˼�f�����A��� ��z".��Ʀ���am���S��<ރ盧���,%��3�t��"'�uf���0UE6��6�;QXa��pG�b�H�.�0�o���0E�+��m��[�w~��7@�����9B�`D��>��F���!a^��Bh��Ů�7\�0�GL��@�Cp�cP�ՒO�"3%���B����Of��*:S2�����V�7�r�����nfҰ�y?�6D�ϘO0G�>A�Tim��l�vs��|]�����9�օ�?)qL冋�3��@�S�o�`u�k+�uo�F�'z�}8�K�q�d�n_|�GO�-J<����a�\�����cR��S	����[u��EI��� �mQ� ��T�k��mGs��a�N4+v�4�|kE���b����]�hm���eHI����d���!r�$j����a�!�E��t�(ZcT�"�3La��@;�n�bX��� ����LL$1�^�Cs4R��H�d4�< �Ԟ��A��ٱ�P�?OUU��F�o�,�j&	�����.:[�mc5\%ߧV)R�Γd�~���d/�(@�_�!|*�Q���Qd	������@� +�.q%$�ّ��]��+�w=V[vG%�O��?r4U�P'��&'�6� ���,� �ѝn�$$����Oo�X��-����&{�WN�kr�Q�̤{&=�n9n�a�
��&����-��{%�W EU='el�-c|E"��aO$��ԉ�Q]o�N�� "G�����u��ۥ��i���?�z&Twנ�V51�[�$���ےtelr�����^�b��3I�ωc2s� ���>�/��_Yt����
%�}�;G1�9ҋ�j��m�'�a��u-maY���)��J��	������w_>f��j30)�Ѧ `��#�,eo�MM���G`���w��2�}$$�F�R��{�������^o��6�v2��. ZpE��g^�6�Ɲ��7�ȦӾ�f�PlzH��V6��@�ߍF�!9����"�ռh��j(�ɷ������2
A����켊��z�	�iG��S�A��h�\�D��j �n�~K�>�ߋ������=����5FdP�8�|�~�`��Gws���4;�?��2��(]M~y�9��2d�����I��82�_y�n�&b:���M��D=�^6�l<UE���]�mZ}|+�Npl��$C,���������薤���Y�]��&��q1��|����O6������JR
��l�Ĉ��q? ��8=�	$?�((B=@�Z6n�G�|d�
�� �����'b9���z��8:�ʩЖ�<
��c��$ �,�s���J�p����ֲ���߿�>�7�U����L����h��.yjr��&,����(��}I�E��[�&Q��}i���
a�"T�lE�$��w�2��~��]5I��'B>}�O�x��B�l�$^����==y ���4��Bh�	\^�8�6��Fr7�MI����E\�} ~�c]lh�Ù"���[�UL��g�y��|?�	���O��V����<3��A��H��ke��q�j�td��#�+Vg�(�T����eBQ��|�����`�8cQ��w��It#0�ڧ��J1���t�<?��ܜ!���|V����K3FJ��(��?x�R��_�D&�ť�´�5W6Vc�n�Ebe�0�&I��eh����h�@�������T`��	�1�O9Ao(f��/J?1;��ͮ�<sA0;V&v�V�k�J�X]a$��4�5`=o.�Z���)a�����q����ȇ�ڞ
�,n?���Y�41�\t���HtE��RIVj���p���pMp0����*w�Άb��J��M>��z;�9��4��߄�3�̓��o��d��]�~7T�����p&�%�B��kbH)�ᾖ��	����ȡR;�8b��u(Ј��Z�-��[��%]��5C�"���6���G<���+
U���]��WD��ֵ�A\�д7�����3�D%�r���>��nҼOFɅs�����R+wm��k��nӵ������\���\�ۅﭤg�����ƃ�.�K>�^��������81PB��Y�;��7��cCq��2H�{IcXL{v��\���H �_Ś(3>�^\�^A��{�jrə	LOAL��1� .+�R��y'����{2����Ȅra����4㯴�����@\�f�o�D�M����$~,�H���~�M�JLn��ԨH{d��4r�V�},�Y!��7*�4���#9|Y�S������m��\��ݩ��S����>%C���{�n1i}1rlSh��6�Ļ��Fh����h���h�B���5BN�%�FZ��G�=�契�a��� �{h该F�G�=	��ܩ�i���~����`.`����	 ��&5V)���ow�������k�3�qD��~�F�,o>{D�4�5qp_���%�!zBa��14���M����i��@}u��������٦Q5(��M�%���0����Pg�L2��:*X+�I]`qo9=[�i!�R}dkDxq���K���_�=-�}�p����NB?�4ܽx�DZ4��)��0�x\��0��E�׋d(^�x� �-5.r;3��}	/�8�\�@�����Ģ��6uKzY�K��4��U==;:8���2\��LJy7��<|?�Q|-pb���Ĥ��6z��*(X��a*e"��xY�@��f��ѥ���6�ČM���AK�Žz:^������� \ɽ y�0:�h����EmY~h�&�l�i�[�DM{����̀�NGǢSeI����T��3��6Q�'�-ɽ��X�dm�vK��@Eo�'x|�74:B��s�QQ3�����Z���F����#�]O����3��{�m��Fp�����#h�/���"y;&�J� �*�P��J|�s����bq%e_��HOW\�!تhѲ$��sh�V��S�l$J)���';�R>�f_�b���h�j����{y3TĞ0H5�uYD�P��BgQ@2�8X�kx�ѫѶ>zf�y�LiZ�[
>g�����	N���o��_q ,��ݜ�c��+�&1@c����9�����%��5L��L�ט��ܬ������Z|Ϟ#��-z��U6�9a|�nSv6�X�L��U��D}$�O$M�a ş�{�͊��\n��tȚPωf�<�?����[T�2����v�5���8��>�D��}�᪝VDr1!���#H3�s)�)���a�Z�d��$	"_&�i�5�d�e����F�c�uG���E"ƚt�AB�R�Z��gC�z�'r�4�z�6n�x:�{|�4�1.��뫆��ަ�N�]���W���B[D�D����#�(�����.-)�5ю�δ�g����i��B�GPx�2��Lǹ�o3��{,B���&�5�w�E�ո���z� L�嫣����>�^ו���J�./��|�
�_~T��A�Fنo���@���Yb�M�%���G�l[�{�%��;��c�I*��l����۴.��0��`�D�3)
p����g6�ф���R9����H<�oh4`���-g���Qؿ�����K0?�:7�ko�㷥�A͵E�A�&�G�5	X�Ƀ�z>],ۇa��߄7���׼#�-h����!�ȁ�J��7�6~�]�Ԧ_��7ޓ��\�ՆQ՟�3QvQ�}>��:.a{UY�4N��bc��Q��I���u5 2%[�e*�N���^���x��4��6��9�g0�FR�zr[�H���zP4�iMk�!0���z��Uo:�F�|�>՘��LۧOzz�T �F
Z1�E�)�Q(&��{�o�� �S�dX�pܛ��Ţ[p��m��csw�瘜@EMր���Q4�9��.��9���9c���x*��S��� VY��Қh��?�M@��>�ߓ/� ���R]�ݸ��qT?H����`��A'���+*d�4��7����/�{�k��	۬t}�i����m?$��)y��O�Ԙݷ��Q9h劆pu#L�%�t @��k���V:�]�*���͕�R��S�S�����䔍�$����q�V��!��v� �Cꆆ���<8�[��x
��VςY�N�燹�<9�/���X��,��������uK{��TL7Z�yN���S�1�
Ŕ���9^��o�e2��/^z¨�=Ci�����`s_z�G ��L��u��J[��*�Z�u-�6 a�E�w.��;� 8Ӕ��d+����bɳ�?���%�A~>�BO�f_����2ʠW7�59�]"v
4mt���,�B<]=R�t)�=E�j9�dZ�)7���C�W,
5�4�����J�FX���5�f��9�qN��Z\�� ��П"{< ����t��A	�I[��0�������Az2����s�0�����!q�xx2ς�q�F�N�F���R��$��P��tɯ����7��F�{�0Q:9p���!�K-Vd��C|TGR� �k����o~녵��9�p�%���CZ�z�  }q���&.���<8�u;�
�'^�H���#�ﹾ�Ų��&[�f8!��B�����ߛ�VQ݌���k����IU f������nN+;��+���?�S,u4발��{z�[�y)�"aD�)K��5w��u�wB O�#z���8����~�L�:̅���3��8
g2"��8�ΰ��	GΤ��f�!�IJo�J��Ȼ��e�r��쇯��,��"��?�yI�Dj�^߰)�Xl���!���G!|�	N�`te�q#��_e�sΡ��pS��2%V�lS��&��޴)�
ޚ��o_����!Z~���"���e/m"�YL���+,D�dhr��C��H���Q�S�4v���ٓ/�O�~<�z�3c-%41\��.t��x�7��b���֥���da��''�7dH%03h��Ó�pz�_�NW@�&��«��C�+�>2�i��U�1�W���~`�w���w~�e@�u�>9_�dA�\�^5�&ϑ�#����9�܃��&�lK�a��F`813���nD������%�_��<��[��^]�\�|b7��'��&��!W�N\������\���stj�d�D�Gr��ь+S���;fY0v,�c�0E��z�@wD,	�����8��~n��i��.�D[�E��z��չng��U�>MO{�� ��#�����gQ�8㿕41o \��R�>j�R��αQބ�-�Ea��V�S��}��v�!%n�,�|�!�Z�5ܩ������%G)���8���<�]FC;~��,(�;�ӂ��.s� +�8[��م�%������CvB�a]#n���i�!Lɭa!���kґ(�/���L*^�WK�[��m�v����@�+�����\�ZM�3f��<Ҫ�E�=��d4wÅ��(g��2\�E�c�w���˂�8���!	䱒|	��̽�w>��������G�Rϥ]�}�+P�8fpDx��M�
T�
c�o)�E5_'�O�y-#��������K:%��I������r�$�äb�)��@� �u��E<�����*�����I�~E���8y;��O_צɶ:����X|��PǠ�iۘ����쮙�P�T�ٍ�uz�cN��p0Ǌ��>q�+<��I?2�qC^ᜱ�t84fֆ'8̞�W�b�x�1ًI�Y��yv�9���oy����3����U7�zx2���{�,�]�*	�[���/��9�R��<�_Ӥ��j�j�;���K��V>fx�W 7��Í��mx�. =���a.-��"+]�������)��H���2���;e���h� ��CTi�_T+�+�nq�H�)�c��S4�_H�,ǻ��;`�hooك�!���/�O��u3c^���0;B�#!��c���Q�#~E�(�O�;ow��{l�y�U#����W�4K��e�O�j0�4GO-s�d�\>��=����[Poɕ���_�
��	�- .��z��HZ%�����ӑ�LO^n�����);Sh3i�4�|�^�~Lі��&"��c/��i&�Lv�G�I>"�(��Թ��L�q0~�h�$���;^�[� �N��h|��c� �ƅrƠ�R���������⨙����R�Ƕ�Wg>^����T:R�>� 7�D5�E
����Z�J~Y�(R��k�+�B	�o��������JD��F���&u3��|r��X��q�a33Ч`!=e��F�Lg��_��j�q�A��r�G�e[�5l�S~���#;������!~s5����R�t��I�Kn��� M�>�?^G=+�?�F��mh�a)�_bnz���h�=7� �!�D����I����2�M��P7�N��+�Z�ɔ���5ha�y撑؋��Z��ml˨�'KS��p��mF(�����O~l��FS4��vK)�D2��b��c�Q�U�L�v
Mr.O|��F�?ǜ������r��]Q�F"�Y����D$6-��! <}f��z��C����;%k^���HU6+��!��%.����TJ�N�]������Bk��J�ݺ��guo���!�c׶���c�LJŵ�������)O��_�Mh�"2�n�.��N��H:��U��r���-o��߉���#��o+G�Z�4�@lZ�&.�G��ГMÅ��8��G��O���[qW9֘l���a�5�p'��3̞���Z ��z�"�"lW��s��s�᳃�|���&t����|�dw+�s�7?����BQYZ�P����g�R��U01�!�a���_h��Ǽ=�R'c/�C��s��RvQկ��"a/X/a�
XI��w�s#8��L=c�b!oLB�^����u�-����l %����o�����&�P�{���d�|<g��B\���G���:=&��+
�(�jO1Gae�=��	^�h�'io�:[r�R{�:�Ydj�x��z3'�z1Yu�b)�|�)r���A�9R�ؚ�L���5�'�zy�Y�����Jo#�����������6�^,i|ZFl^C�&���ti���K$��������_�O�[]���u�zW[��j)fv�KɂQ'�z	/ͅ6k�^<:�����m)	�,~�"���~��0K{�W񇤞c%G�9�#L�Vӕ���$�pLx+?&�!BeP�b��v����H�X���G!�֢v�ܳ����o[:y�Q��R�
� �;e7r�S�T��-X�T�8��d
�4�Y2`l�'��i[(�6f�[�2�����v�a�4��*���uQ�K��bMe\PʪD�7C�� �7�=YI9��5O6��ת� z%�;w��KΫ���c=��D8���>J@(^6�����--Ka8�&t�W��=t[iG���|+�C?]��E9��W��I{�{�MW%���{"�I`�O��%����ն���C�/�7���"I��(��	��2A�`uE���a�Z�K��2��Q-��#+�{lp�u�f	�6�4��3k�ZT�r*���GNE"�"lZA�s��'�=6�2��P9Cʈ�]��g��R ʫ��t�7�Y���k���"�f
�p��[D��s φ�{%\:�B�ͯ>��	�5��m+��ZH���R#o�B��rCo1}qt<��-�������̃���E�������Ҟ�����RO�����^XtGRPjS�qP���Z��t80�T1
١H��^K��ՒvY�� v��D<jv�m���.��\	�A��麛�ya��D.$P�g�Z�ҟ��͟0T㦶�A~��:-�h����#�m�[#��y
�Ӧ\�x�_(�{<���jx+��h���2w0���.+�~���&�m[�쓺K5��NxI���:2܌Za���{��F@I����5�<��X�X�Dng)w�r�^	��k���xl��PP��ĕJI��g��cC}dcx#�P�~1,+0_��F��I��:��8�&l�mʧ����+��b!��\{�W�A3�Ae��S��n���'u���)>�� hW��-��K^M \f�a�a��q~I�0�kw���cWGv�ǯR2��:OE��dj��F�ĭ�yZ���m7�0/�~N}�F���P~Z����!e����4��I6�F�݅^{_=G-:>d�Pt��w���1��yK�-BX]�X��� �d%v<B��H�Q+Nh4Cc4�h����
����c���d��hI�'��ĶSv�/��m��i.��F�0��C���+��M5���Dh��\�v��9L�4�>�:�5�&�0�|xZ��X�po}������h��y��{rb�����I����k-KsѼT����|�ok;�hC_"���f�H�HK`J���y�|Y��'���
�.R�i�P��ol'b����QZs�t���ك0s{� F���İ�u3��9g[��b��_8v9�!��D�=q��`���+fHNFpȤu��@�D`Z�ט��,�Gu�i�A��_� :��7��t\m��[�ׂ��c��2���E��	Xz���<�y��'��~�j���C�������2AۑÚ���!�GtG._�٠)L_�y��#m�O��T!��o�ɠ�L�H��3���HK� �����S8L�U~�� D�z�E{����*�Έ��br�.�\�a�,h�X���	����4��}A-Vk����E�,�h��۱׷�L�3<�*_t�˘'�R�p����I��%_*᝗G<���"�k!�0^���gW:YC��.�7JU��v�l�/��8�^��uMt�|����|�j��g��;�<�r�J����y��O���Y��36����G���M���܂������O5˿��,m�����\`���C%OȻ+T8��ui5���,K�K�P7�$�0Ɨ�Qt Ƹ�+N�H+���#@]�oG��گ5<L-�H���� :)~wj�Y�Ecz]q���Z���z�{�A/<"I��p<�r>��6�,,����)B)mbFH����^RI}��'>$�8�~���@Z>���-��%���X��k.�H�^��[�l'� .�K�TȈh���i< Gq���za����Hd����4v��K�.ſ� r*�#p��ru�d�%�ҩ{�m�����x�ņ�lZ9��"&%��.���,I�VجI���s��~�p#��>5do�[,#	�"�ba�~���ƔP�%�,:]�*�����J�@���ylN��$ ��޶4O�:��9b����r}'�s����V.{��²ف��S���C		������ ��iD�����M�5��H4����mŭ�BO���$�E|d�-�p�Ɛ�~��;#����󟅕��DCn`�j�s�B@eX�δ# �8�I^���vP���)-��ɰe��OF�[d�v�A*ꏾlV�ihw���װ7'+B���3�X�Z�[��ڵ�A��t�DAH��
"#�e��$LB}ܕX��#d�">�H'n�������#+2�ѽdj$�3°��ݶE�^ГXr��/K%�Q�oj+�h�!m��dC��2�3�������7ץTT�VO҆:qS�AК��智�E�n� �X���@(z��{G��N\ݾ:��N]�7@��x(u^:f�{a���`ƆF���Ch0��P:`D���^�g��dW/it�"�/�\�$d�1Q� ۟�,���<��vQ���Q�[[�	Q�2(P�N��F
���ۿ����y�린Njk/����!E��'����>�֯%�lp���w�9X,G�jr�%�f�,/����k��OѭPFj��!�w7Dݣ�A��d�������I9v\L��wˍ��� ؊Ury�p$9����4 ZL�,��5�q��׌]4��2G[��R��U�Z��D'�"�I��qS����2Wj6���nX�nC�b}A;�湲P����!�$�g���~U��μ�jC��퓶�~�����+�rc�
l��s��$�.��w��wJ�B�pƧ�'F'�B49t���ۆ��A��'Rj��+JQ�2� d�����

j$*�E9ٝ2���x26yl�,���13Q���R"� Mn��^����H-�>�6l�d�W���^rM��7��ϑ���A��&f�y	,�B�.����X���K�zs������\���tǏ�oW����%x�7�%�V��p�E@؅傛�bf�	��@#��hT97I�b9��Ou���"��B�I�#�,�U{�����Y��>��S�#;{���,�'�;\Hz^�\��u���d�vq���>�s[���k��g�.�UҎ"a��ZՋJ�&���٭������d��z
{�^Eն�A}2`d\�4(����.^C6Ν����ͧ=/�H��!� �O���֫_���gA��hy;�HM��Z:�Sb�M�ˇ���~��"��>?�p�+{�Nhx�Ѓy��f���?��Qĥ�\���J�J����o�i����+s��UvH�t5�:&A�#p(�ι���:���Q��Y�U=�>f�6�~�MF��6yW8�et��T�+@�?����˯H������o)�._�H�P��6�|d;�pϒ��:���,��9���`���p�l@��r2,ĉ���)�tj��ia�&�ڍ	J����^<����T��R|���9q^m�d	�.���s��w�L1qr.���^��������^�����|�q�-�.SS��6��ʕ_�9�L�I/�nk͌�����2�D�C��>)8��_DC��_	�[��"u����I�����*��hRRn��E4�l���<i3$�ha�H�*�MO�ɕ���Y��,�D~��97dT�p��UKD]t�o�N?��էC��G%P`��=m}���M��r��+#��,	c��HۇtA��6�ȹQ���᝺�tC
��l=~׽�B�2��`��a�/�O�>����2�����QA��WЦ�%�3x��?%�I(��u]�_��Xk��co�W��)��\�e��d�4�ч��oGU�X/
�0������'�y�T�h�&�qvX냎�f�LN3]���v*@�%�W`�Q(T�AU�����Y�	��������b���E�?_t3{@�	�o��.(����	��{fj�)S|ָ��oz9�^-��#ύ-�DJ�N�7"M��D�PV�ﵮF��b�~I�R�7������S����gӵ]�7�]C=}�.����A)��G��K6��n}���D����s(PY��½�(f�M��2#���Vj��*�WIR�����#f-�`t&B?��y2i�N6Lc�I[�*�(!�%��Q�ܜޝ���"0}�;�pmc_�?�}.�[^	��T5��H�%�;L���&���;>�qQ�K숍��΀��Т&��_0�ĺ��-�5��d�a�X�č�;L�1��}�D���}�r��3�3`=:g�:��x�[��?�1 �7�O�7ǉwe\�p��y�(Г�̰²Ǚ\f6}��d��da*;��t�)�:�Z��h�幝h�$n��0J\vn��b�#}<R{���ל��=5)o��f��t����Er���_W�ݤ����LS��ySPe��W�����e\�e��d̉L�=���tJRbQO�Q��ww����]4�p�X�|�خ��xdߔ8����&�I�"�n��M�錢��X�k���� ���0��h�tFgP�MS�,���b���¡�񶀩��S��E+8i�Ri2J)�q$P���1ҕ5����b���e��YbTEnW1Ω20��w�J��6�퟊��HgY��1fLt�����M;�"F9��=?2X�T��`;� �_����H�� ����d���Sg������*����ɽH��]��ud�`�;�j8�� ��1��U�3�xL0�����m����gc&�eC��zOM +�N��Y;E��Qr!�A�$h�kG�$���FੑP�NHh�͍ܽ2��<����~��L��p�!���I|����:F=r$
�h�q� �?L.aK���ڃ�ڒ��������Lr[�X���^�~w2�.�?;^(��ܭ�P��| MzSl�,�A��ʾ�"���J~1������`��E�~$�)��:�7Yq�£�e���{,�R,6v���B�nv��v�V��F2q�SI5Ȭ�K3*A��:a��SG��h�] *�@7e�����D��+<�nˊ�9`�#�a��_� \ָ��4δ������9r��V�Ú$�(����G4D{ʭ<x,�vA'S�<BP��|��!oՐA���-�x��9���[��"ipQ�)��� ��}#}��Z$�ehVU���B�_QB�q�Z�f�'l�x���t��4��ļ�t� ���7]�����S�o�)��3���Fl!C����G����X����&�� f�w��g| ��q@��sW΋��?`$�~���5��(7���mQ(fnA����܏�+��K�wr<�\��q��S�~�"�t�N�Vh�HJ���(G��Ml�?�9)�a?��z{�0��IգIU@�|fӬb�-�ѻW�Y���b����l3�����ŉy���Iq4'-oE��P����f[��lH�;�l?��p��"wtuCs�l��չF'���>���t�ώMC��5;�k��Q`�f,-�W�V�G��W��1#�ueĂFdmg��ږ��3Űn��bI��)��O��-���	C�7��������%�0d�R�{� -�Ј�ƚ�$�{ѝ��Ǔ��ߊ~}������m���*1u��"��u36���5��z�>8��,ZЎ��C�>A}"|O��|H�;#��(F"��_��m���6cm)<���<gk��TAJ����?���&�. �5~9?�<���#������)��{vTv��,�N 9`0����ݕM�z�ւխz�ڱ����7/лULL���B� ����y�=} 8i2�5�F��%~�z��I�#]d�C�\F���K��I�h�~K
dh����^CT_�b�~��ŋ'�<�{��ew7�&�^r��1�+��Q�5^t��&W�oB v�`��b��>�<d�Q�8f�+f#? Ȣ]�TC�fm�:1�"�1�B�>k���J�VcUH����X��0^E�	W�]��X�U�Q`�B�*L�O�*�ʃk�ݛ��o[���b�gr�`�c(�ޯ5�M�.ŕJ��Xj����_ 2�rF�^�8�m$B�l���Wj�-�Ha��Mft ?rC�{[�g:k�3�"�{>]�@W1��@��"�G��_��h��l`�+P<���M{j�I�]HH���ž�1��a���N��Xh���).�Ô���韛�;���L��8��b�]h��'��L�jn�O�#f�uKh϶��e �D�꟒,4/J�W��t��5+���8Bb���Um�0`� �i2��{>gvO,}W'S���% <�,<�Ef[|iꗕ~�SshW̮!>O���4�3������Hd��ˎBd��7�#�oJ~����h�RCV�`+��K��i.�v0�34�RP5T��7蟸[;�y�VdwIj��l�K`�S�j�(Z�x#�kJ?��Κ}�Rk�{�xh]_�ҹ��	������ث���P�v��4.�,u7���玡a6��M͜F�n�0����$Uk�ȇ�I:�`��p�L9���h���aG�ᣦ���h˚�Y���D5xe1E�w��R�����5F~$�Y�_Ҹ��KwI��V�u��L���g{��r��﷔���#�W�i���JMR��i��|�d3 �^�,�������$q)�\ LKxq��,-�&-��5��Z��܄!� �)A��H�Mz�z�,���.��{����8;.��G)� =r�FI�bǸ`�<�j����k��++�^?��P��J�P�K����n�kzA@����܃�iMQu�>�MT9���s!=���B����1N��Wg�޴����+ @%\Y�|�b�����a�d�I���Vnr�d�u�uy��P  V�NU��Ȍ*�0���""i3۽0:KT��tEw��F�^7�~ƛ^H�M�{߄x �$������.�����4��fI�����w���W|3Ԕ �H�z&�'	���;��ғ��b����m���8ĵ's8U??���Э��?v��(������Jhp0��/�^���%*'�;��?���ԩ�@%��K;��p��F#dG�?M�3�G���s��j�yï�g�T򤋤l�Sj�c�wpD�6�C_����D��+��4l���� ��ɫ� �M�^��<Tۍ�E ѡ^����H�$_���t���\��yq�~�an����x�:C>I��@��5%8����l���o�}9��ԫ��?�<��h������7�,'=�����#�"@��M"��r-*3��I���)ޫ��}�4�~gP��+�f� ��6�Ĕ�#3R��
C nd��I(�m q&�>�r}o,)��Fk�VU���%�S�cT=��T�>����I�7�6kH#��q�߮Z�-�����y�rj���|*,C'l(���&��h�ף�����[^�i6�>��s[�9�g���{g����D�����ފlj�����A��̀���X���A��h�12c��xoNv��>\@�+�>��ϫ��CVC��9c��u�DR5rP����r9������!��ÒEKV_���}�%6��]�(�����Ğ~���L���U�l�=�*�����{[�Ԇ�����uF�
W��J����r\e�*�|���@X�r���6�Kp����A��'�	�A"��C��З�������0�t,�k(I���	�j���Q���|�y���`O�/����[.�F��Vm�e6E5��1��.}�P 2t�9�t�y*t_!�'�����qJ0ث'��X{���#'t��c���U�ny�7nwӚ`��D�f�܈?A��Ȱ6��9�� �|��J#� .�4��(7��&��M�8��*�:�IG�I��t3Λ���	�<h�7Y�Q���+%�aЩ0j��_��g�X�u`�MK2��+�r��Fid�Pw�������H���>.��J�"��_�/iMX[����U��X*����緍�8�c� �Μ�f�W�3`n~ĲHO��ݗ]��x*�!/�i���HI�O;<:0������51JNL^0��R��Ф����ZQjV��n����SN`�Mw�:�����Ápk7����Z�m���I��\��P4�0`�C���ZA��wf��l�#�V��r>]
�Jl�R�ҜM���[8wT��,��D�znT�g����g�+�#�����l-���e��\j�ꆍĚ}�N��;}����?^�s~���.��xZ)]X�`�����d����ӡp�!�B�t֚s��UC�-NA�=�VRN~����>aޓ��W��>~�B��JR,�U0�T����vk��}���\�_��
��3ҳ�E���z�W[de�L�h9��t�V�l�fc/Y)J���'��h|=�S�ݽ�SZ�|��,U5�A�c��Auz�K���4�[v_�ڴQڀ�.�0/�;$�r�4�^�lR@��9*j�E���v)���J���`d�q�V^�Rh��]��FF4��#i������SA@A��PGu%^f����Fl��+:���p��Rg�|SY:�)��Ž�n�v�1�GaL(�������h�輧�<>��������5�)1�S)�T�-�a�X��ꢓ�Ѡ5%̉�0��*� ���'�&0x�4����x_��|��0	�Uw�j����R��ԕh@w�1{CO�	�c�pu+�=�瑟�� �"�_���8�m%R�Z�_W�b�Fr=��by�l�R��>3�T��j�Lm^>�[
l���)���:��'F�1q����dTڂz��9�jݫ#:���g�w-�Q����ʀ�X���ޮ#+�RGײ��X)v�{R��WD����@������64C�	��<`ç���t}�}��*~���G��:p��Į��_�
+L�R0��ba�ȷ`%[j�Y�uD�������hܞ*) COѨ<":�=��u�����Ý�i��&X�7=d��%��r��/���Iq�dfO"���Q�}��t�;W%k��n����<�dO��E��}�rVJ�����It䓢J�GO������GF�~��Z�S��'I!n͆>XU�m��>/,O3�i�fZZo�Uj!��cr�լj���>&uDYd�R��� l���)�əZg|������� 8�=&U��P����'#�B8UO``2��q�Gեo�F3��ɩ�C�VE�+�R�ҹV�e3G:��u��fkxnG_ys���֕�^[+�E�U)���O �<��2�Xh� �[ހ���Tc�L��_���1��=�K��f���7
��]u��[͠��H9��k`�<�:|���^?s��k�+�L�l��\���']�d�����?��Lr��B;}b�Xm�	m/ePJH���<��R��ս�y�/��	!Q�&fY�
���6����Y��ҟlRC�y�y�����wI�;�����U�sҬ���wRҥ�g�;i� J�^#~?�����JK�3�R���O
����5�������޽�;�8��~1�%��N�]	ֻ���n���~fCR����s!��pܻ'��p|����\ȓ��(L[z�ĵ�i\eh��iE',����Ȑc��/��dɰ���q��ȝ����cFE3���c��L'�e�A!-�1d���38��� W�*�l<}�i���e��ĸT������G	���bW�e���5�16��$?�᷂#�-}��ݹ?x�_��fJ�#�F�$����N���7Z
<r�s�]��rS'�!�9HQ ���Z2��^ںBfl������<N��D����32�БB�����5$3�p&�xA	շ�EO�`?�`p��4h�0��~�FKisD<��UVߔM�|�ԛ��@Fw��5~��M�����ަ?�w���	Y����li�Z	��sD�'�n�
XM���(Qy7�0	j��I��u�������U���.���U�����z��'��H����6]ڔ�PE������I{)�g�V[����L�?���P�+?8�RE�׋�f2f�7���S)���H$	?Ul�gĻ�^�]N6 ˲��9�a�Ǧ�I.WN��ԥCjy=�
e� ��M�*}��������P ���[6{�k�
��u�'.�Ȩ'��i��:ף��|Y��%�^�K�F㍰��o��4��k�~��u�GVNj�*�����oVZjk{��@4?���e�	�~1Y�E���	�O�����C�D_P�vU�gyjڍ� ]v#h/@�~���f��U~��_OB��
� �E�m�u�o��Z�D�Th�!;i��{��>��o]����G���.9�y!�b�ص�"IR��;s���f�$�,Hxe_4�5<��������?�u�,)b��N�e;Vأ��
�;�L�8r�/�[��
��ނ/�b����4�`�[����Q�u�W�Y���ˆ�zm&�O_�Ǜ��3ڿ]��L�\,5sX�-S�ܙ|�����ĮFFɼ�����x8�	������ׯ��>	�(͸�q` �o�@��*�����t!��>�u�x2��d��\3k�ORGC�}�w��>�S>X��n�$j��u%��'�-(��D~����~���u&�6�ծ��
pƠyr�[�s�,U�j mֳ�6����Z�12��������Ky��ȉ�K�����$-ݺU�4<l��ꑦ�{%jo=�o�����6�!j�i'o~�m2�%u�e�Qy�-��d�I$���D��.��׿��WOX�� }���p�}��5�Q��T��q1Z@qaZ��Y~��z���q�X<Cr��j91��ʖ�5���'n��o햂G�� v��φ�=�(���W�:zE�k��JPe��G1Y�eX��A����y�muZb��}�~����ɀ�2w���0�tb}�?���k��ã��k�}ȃ�t]<-�~#��x��0q�}�*��)^!�"�u�B�M�t�Q�U��H�~σ�5<64���s>6�R�˘6(��B�Q
�6RW��oGtj��ԭ�)�:|��X^kx�Fq��6��_fw������F	.D��._���-܄ߢ8iiZ�ڰ�s���'a�m]0tp�@�Ċ���j��O�=9��q�V-<�K�,�W-��QP8{�Ԥ��T�&��um[[F�Ն7�ZQ�s�mQ31a��/e3���(�����;3�+���_�maf������8��R�{�9)�Y�cp�fѝ��yɍ�P}��%��XP_<��0�V�J(b�����RL��2ב�qؤ3�'���D�����i�'���>lGÉ�s|�����
l�vs2����7	[���ݡ�G�*�zU�\�8�T{F�]�V��T���� LL���x8�$ފx�{z�9�7'3����e��v�W�W�n�6�l������W�@�zbE�`���0 �v,��cg+���*���K��#{�Mֺ�bM~מš��������sW��3Sg�%w�@���@��F���e����M����SA�<�N�>��*X�X�1E�����"������+�e���G�����l �wOſ5�/F-WK�ʕZ,k���7��<��s���_"�>�1�e�D�)������L�6t�:��<��%¦��f���?����5ے�C�d=��y��o3�a%�	��D��+�Z�q-�*:~Ȼ~X�C�Rǖ%pa�A�ߋ�F�K�.�_��(a�׋5�1�&qh�����|�ù�}��I��>�D	Z���''@%����P�ӥj�7�.0�.h�ޤ̾�s�
����{u��zJW�9{�0�����SM%�Kr&��
��-(ha�:i�h�H�!���yh����*r�+l,��Vc��SJh"{/�-�W3����l?*s�w\�XB��z�jG�Ӫ��WV�[�b�����Fםz�HEj5�D��zـ=ڛ�W�.L��}�m�[��d�A����Q&��^�5�S�6�+�z͕1���8~^z1X��~X�S�x�+�Nrg�A]Թ,[Y{ds�>r3��f�'��r˟*�k�I؃S�'����q�6^�^�]8��n��󘖪S+	��wa������ڗl�A�O�NHپ@�'�-�VX��e"�
(ȋ&z�w��$dC�O��n�:l�<��h���Y6T&���UF��S�U�����$�0ssQc,z�ҩ���^��Ò���Q�؁���ME�p���}1��{Tx�8�ꓞ����AY����p$���'���ՙ|鈥��W.K� �T�x��s=Ţ�Z���q��+ݟ��`h����g,��ͳ�Q�=3�կBn�M�O.��s�>��Pv���]4� ����5���dc<�a���ؾ�����3~���l/���,\�CO��\-D��j(~d��.��q��t�S򶜞:ʧ�+Bg��Ƕ)��B��W�`]��!��d�m4F�H�u��@��_<���`R��E�<�@�l�eL��ߺ�s|+�GA%�/+���tcD�9�Hj�Hn���ɜ~|�lm>N������3L����
+F��2��,Hp(�/#�r���fV�+}�+^���#?��բ��y1$2�	���R����
Qֺ \�je	�Ӎ��H��d�yb/����mR 2���,��?�TJw�]U��WU�D��t�RO���wM��2e�A��[��dzVw�W�����4�3��_�_��a(|�A+ʌW�UA�u�A�;��A[�\����_���lw��r0t<{TVL�x%k�,�}��������`�6��Z�77�¨�j����5�LM�e;�Za��1P��Ur��^����dx4��3K�n
tꌸ��B`M8�gq�wmk
ے��ct?�0�q�&1���5���8��_�]�MJ�m�f���h��WE����c��k1�E�K�읹z�f��I�#��n�ו�S�u}��.��4U�,&S����C�Q1�����7_+><5��¯���&ĝ���: X�S�hs�踰�����,8�Aӝq}�q�&s�N=��e��,2]���e�VF��4����P���S�2���-�$|YDm5����4<���U�I�tl�!#qqI�������Q��M��#�$�~���x��o�8���a���g�}������*���#�
�o\fh!P�q��%6b�Fq� �O0!�e�?�U�dX�[�=�g�6��KUᘤ�����V=g��2qS���f�E���Ƞ��J?@v�et*R����}~>��4nG�n��!�O��2i��h�v�o��]��F�*�T�)�ݡ�?Կ���w�����fh.���)j����pZT���>,|^BO�.%nV��aC�7������=>+ҥ<x��N*�1l��gC~��WJ ���w(<��H`�^�C+y��$���Cq:�3"/��=J��t�"o��kk��(�EbѥTFCM�5�;��DB"��؁\
n~ �+DK��i6�^]�1y�jh3jE���!H2K��F���N�}�<��/x8+s���`Kޖ�ׂ�\�h[}��xw�oI՚��"�Ֆ�u��n�m� �hL�[H�=ω�L��1`,�\�j.�l��^���z�j��u5q�&������"o�����<����&!ص�2��ۏR_���\J4Qa�E�=����L	t������G�kj*	�m�F����x;�SX��E{���
S�ʩu��>���+W�m�oK	���J�vZ'�
d�NP���_�sDHQ�4�T�Q��5�VBy�9�k���Ƶ�f�4=<5Tȋ2��.�t[/ZnXUP ��
?��� �(��*�0���v�Ѧ�5{���l��G���	� ���?�����5���J�*Ϋ~����ޫ�^S�4����~��$�����	�)L~(.��Ѝ��˦���v_��o�V����dH[?�
i�WY��}[R�]bp���ߎ8i�ƫM��q��������z�+����V�X24�s�"��iA��~�/�Ӱ�^JYO0Ϋ���{e�1�(q�g��-�v �|�8�ޣ�� ����"����MB�>+`�2-<��O崦W�Uxpαe�JM���<��IS�㈗���O ����}*3���w��)�ƣY�;����ْ��ϨԆ3��@&��^X����<����O��)��K$%�����ڀ�Ռ��
�Bg)��	�!��k���6/��_�X��ư�+e�1{\�N����d�cYЌm&�m
E��L���W������-v,M_�}�k����R<�K�����YS�<R~���k���&,��t[���8FQ��Īނ�F�Ž�y�o�3�|��ҲL��}YS18�6*��{k����j�Q����l��Y<�/+�M�/��p�y�CU>���SA|^Ll��G�n�P�?2m�GM��BzI�$I�`�u�KB9[ͺ*]n���{�ֵXI��Jj��;����u�>n����hN	R��Iw[���TKf���"(!�;�f�ޤq�����X4�&N����>����m��>w*o�'!
(�a}Zd��tZ�@6����0��ߪ�tgƲ�"F��"�P�p��GՀ�.>|j�4�jԸ$��[�M< ���-�m��=�} )ۋ�C�cwww�RB�eS���}Ր	k)|y�VA�7�`�1�ʗ���ؿ�
�8�	 g�E�����Æ���d#ӫ�@�!�}l��O�yA�!�ƧC׭�?��;��f�D����U�Hm�R�+�=۳�q�FЌ�Iqb��ʛX�V��R,�9���ǚ��&����6?`G�#�IG~B��$^0R��[~X�K�~�;�(91�'N�Z��^L�n�*�L2�M&��GW�+t��S���_���Ӗ�;L��S��޺�sWN�ӓm�$Xht^(T�-�ZG�H�c�$7$	1Y˫��&>������B���Z�/}1=����l0�A�L��G�|B���uQ�>��CF�[I�WD}	��}7j���y�*��}���O��X9A��4���}z��g���'��jQiy��j��B��pD���:V�>�!!A���x��@w��K����[@3���Wۙ�Qɂ��ˑӋ�-��3ۄ��g'n�0�Pw�:E��yϋ�<k
@;>U����bԱ^����ǥ��?�DwY\��5ꋕ�JD�Ӏ��o��2f�!"C���L������!N�̵���:���=S�6�\j�B� ��v�W������~���*��S�KL�J��,���?���s�59I��q�TD�T>Y3:K��T�D'b�������nK�%�t�|��9��z�p�ֻQ!�(8���RP�����v��p4	C����h �[��-��]k�zXy]1l��eҏwQ(N}�)��͚����H~�u>r*���:}���1�7���2(�h���C{C��.����x�
�Q�l��
x߀�%oƶn��+�ן�̖�(߽�+\��.b�Ҹ AS]�'㹇�+���'m����x�s5���[�U�m�$���h�����Y+��J�JR�������� rP!y���C/�g�*zc�`���Ө��]��!����3�`��_}�O��堁��R~N;�ߔ����l!׮�m��g�z� �]�1r��US��h�&'\�*O{�03�Z�1V�9���3PgM�����q��@|&��!M�;�6�
� Q�w1��)�p� (�ö�)�)LS�Uæ�t3�.���aDn��|��Iu�#�_���Q�7��e�M��p6��j4��z\����M�R}�p��'�o1G<]I�M�>�^�t��cH�mN,�ķ���l�0٥�8Z(�</[F&h�;Co���e@)��u�U����?�$��QBf�F�YU��4ލʹ�ZND���yu�Rw�-�d��؇?y��o:�7������5��q��!K�����8�Or�#�~��]�6!3ܗ�n����y)�T
	9�х����O�@d5��6vp��@sK��J��mg�bX�����p�x�Z�&��b�#�,�Rx���	�M����ks�g�(1�P��NUn�@[,(���{��v�W�M9�����r|S萘(�K�g"t��Fv)�B��M�c�2��R�b𸸴"5� fm��b�Iƿ�j�}C�	�9H��rB�f�8GtS�J�y�z��]\ ���I������]��L��
SP<�Z�r i�bd��@X�����D7#0֋�Y C�R5���$M��Į�=�T��Rm�e{u)��0~sָ`[r`��E�Jn�ᦐl��p�u][ٮiW��S��E�f��zB}dP�:̂b��A�w��)�&���Fc��E�*2P��\4!���x�i{��u�T�.i�����O7S�Lמ1�M�w�JDd�`rV�Og�;E\�����6q�:��;�=M-��.��ʵ�Y�:��Ov�i4�Џ+7H	�;F��h��઺�ɫ�ͽ�ACv�τ�^�&��S����&.=��~,.�%In�� '�gw�vA;����K��mE�UE�,�Y��h�8d�,�_DN�{<�e������f��@�m����
�{o�ShInޏ��Ɨ�3پ�#n(ۓ��d?����x���?��Ӊ�P�"v��K	fu�JSF��}l�j�Rۄ�hx�u2�Ң��|~���E|�P�ٷ�U�7{tU|�W��Z@Gw�<�"�͈�^ԡ��&4t4�Ub�[�g�8)�Gץ�Ј�V-����,"&g�Y��2X<{m����9���.>$��#L��B�G��CG̱4ld��jΩ��#��K�L):�U��Z�i���UT�G{�CBI��G���ک�����X����eI/�2雿��D�yM��[M�U��U�]\yB:��d�9��#�mMCl5(�E��Q�Y���Y�<`���������b�����Tك�ǫ��+}�\z�Q-�XC�9-�o4K@O�~�������#W;�Rc�N֑�⢸huɕD���G�`<�1�0~x����b��r���c��d����s@ք :>����L2ua���Y��<�L��gR������R��JH�a���*N,^�b�����m�.���8�30���I���2�ǳӖ�Ajߏ��5��G5l��_�k�R��YuD,��G�H|�*r;�	�+'zTnxSh
p�񒛉��iː������$u�
�My�A�Kg�0sӇ׮/�~�[Q�>��3`�g��2�lpW�7}O���kR�=$'�w:�����K�>R�������ޑJ��� E�Wo8�zJ?X��
]{T�I�jӝL�#%LEV�Aq��m%��L� �H��0"�'��K@��.������B�+�3n���R��^��^$w�~�U(�����P �Y�w��c�=���@O=����]D��_�}bP$Ү?e�S}�V��Đ樊{6�N/�in�]�У~#��� �o�'����h�-����t�����3Ï��=�9�.����p�ٜ�
pOv)���/]��]�+'Ӽ�f~=��<��@j���]�A���KT�֞?T���*d��v�r��=�.�u�m�����(�10����(���w#�9��B�^�˟U[�:��zn��ƨҸ,����ФK|��-�^pއ��m-�a��,3�h�R�Z�}�WW��O?�_�y�,��t�ܷ�`vh��>�A;��Z�S���R��>[5S�����k`����A��#����P�ݚb���~��M풂����C�\Fͭ�����+-����fl��8�Q<�9x���	y��ճ���g�2�@�a{T/���C������&�e3�9@z��Y��p����47O;��L�r����ld�k���Ѳ{����Fɱ0MZ�{��c�;�YȻD�I��� �oI������c�.����W��y��:F�n�B��}���7v����KCA6�~~�]��	hK���k)����<q�Ը��}\�2C�����m9�h�O
�����m�����%3�2B$���d%�2F&&kh�f�?���N3�[�َI��3#�r`m���FI@$ǡo*%�<��P��%�ِ��N��qh-s\��8��>{��C����>UQeU�0�~>LJ&��9��Ձ�#\�,�l"^/]va���݄��?���FśA���	WKg�~�@ؚ�V�:r�.������d�8�v�Y�0����"�a^��%��7ϻ��R7AC���>nO���ٓwl?k ���ϯ^H ���U\R�8�a�{�whh\��	ț����@�ΛK�a-�<am�9����I�->jIg��!pM&�	hks��9� �J)���Tk�H��7ƒ��z���<N�s~���M�UK2Nk&Jn�<��h޺���?�r��yd� ���9�B�+7����[��Y5����T�?�[�]�U�0w�d$K虥"��o��y!����t|���p*8�}����vf�a�������^M
��O�fy�t�i�̒�����M'����%���etĪkbD�A2AXG R/���C�T9������F��j_��cu˖�Qt��͂^��xC��R�������m���9}��6Tq���*Y6�b�>W��	��V{/N������9U���̒�O�5@��e��c���y��8}��r��'��_�o^��y5ֲE�q�8K[(w�X�Nn&}�g'�v4ݹ���#KL����5o�45�������i�>l��.�GB�@�ǝ���6�U��;m��I[M`)ϱ\�Kw��Nh�!n�Х�%�IF��-�����m�'���E����H,0l��)��#$X�[�j)'����:r��QV�>_4&қ�Uڞu�%m����1j*�w2a�yH����7r����1�5Km¦oݭ{z9��˂2���J$���ie{q�<\a���o���#j�z�뫂(*t�Bl�e4Y�8.>!�!Y���V�uI�GqM!��Fk���V����t��4+���Sc 3��ћN�8p���n�F���;l��f�jl2�&UW��U YV��Ȩ��H�����(C�59>A7G�x��Щ��8�9��W$�5�W�b�0�a��*�?�CҞF��+n�b�?�i�U�¦�
5E� �;�>����1�%7��|s�z�)�V%�~}�b	��C�c8!�O}q}Au���]��N�"��<�|e�{������wm_�k��`�e���m�ЀX�D�m#R�[,9�4L���l����]�����;7�<�&��,*%`��T%��V	~�I��Z���%��:� �i����6D�N���VDM���\`�бDOҩ�����>kT�0�ԈDzz&�{OGIA�U�u���a�g�71����\�cb�75����i�`�9�mig�blcF%͍���CgfE��ͯ3��(<�&\��hp���/Z:#��͔,�� ��f�?�)�/��`%��<l�@|#'Z^e�����확^b6Iq��F���_�:�JC�c���Pऄ!�8�]r���5���H6��{�\��5�=Ě`N�+0��ƽ=E��[�02�lc.=������8���F�A@�*����}8�����d�`�E�.���L>���Ϫ����%.ʰ$��㜍U����H�{~�D�Jћ�SM��g�:��@��S��fRKk�!�^P�4T0�L1�R$h�  �*?�m[���m�Z���n�$1�!��l�0�Tk'�L`ƺ�����t�co9�2�J�9��S��b����ܲ������( 6��i�!�_gOr�]n :t'Jgx$���hT�2N� �Bl�J��8�,�L�@CB[�����BH�E!��?~�Џ��3�Z��$�/��n����Uv���A=*]����'�V\�A����$���:��4շأ�b�؈������0�݃Cun�ă�8�����'#����'�Z�8�%._8n��\�m��iՠy).K��3,IL2")���la�v$PR�������EF���-�xε:���5�to��D�%̸53�J��}�m�/�Q�r�=��
����S�1-�؞�Lϔ�a*�][�s8���p�`E��?N@AkOu��P�$>(��5������H׀�ȏ�<�UW�t0�2�PGF�y��oLx�6�v��U�,	���ث8��Abj֨kS=��۸W�����Xw���$��M7Ar�I�SZ��X	ڂ<7p\�a��P�	�#bk�{�����#�}�W+��6:�{�nn8Iu���9��ڞ+\�8(�.�5цH:8]D}^�F%*�;Ö#E:���%���	��	O�8<��8֠s4cQ y�S���x(�#{��?��K>t)��6� %Ƶ����1���<"�͜�ګm�d�dWҵ��96`��8�e/�#���W��k�&۾��oہ���l����)P�|ضCo��  ��f� ���2y(^e�b�ɾW{�[�"Aħ���5���pѮ(�o�]3�*ė�
����9��)�Gy��&�a٘ :ìB�B�|�	0�aܣ"I��
M���`� �A��"��u}h��;§��Wz��~m�[���w�N,꣌��`V�cS�Ç��=?���9�N�[�͚�ǕajO;w��DuuIIp@E-깗�4��5Dw�����Z��Mkv'!�����alĭĕ� Zؘ'��rd/`5�Z�P7��o�6�?���j�b��Ek*]�f��VۯG�����7�����-�Ȱ�Gvw�k�5��_�x#Z�Pz/��Ԗ��|q�(�gŔ��L{�М�b ��4̖8�3�ʗDeB6�j1��<gw���HO���h`�\�؅��*N��3�黩���׎.x�������8M��mg�t>�S�ABD-т[�=�����au��~�+%t�]16��#��=�%�)m�Y���ė��4�7�s� �����S�PK+���	��������d�r��־P�'|bA�t�s��� �'��x6YR��D���K�|AJ
�X#�t���9k��=
����F+ ����E|�M�k�y��!,Ƃ0!��hA�*)3�Ty8��L��-���y�&'����l4�"���t�^�Oa�;�X��Kq��	����=.L��l��Bu����e{�u���̔���ow����NDҘ�O�2�[��EcPK���yri�\֥�GF ��Z#��N�C�D��VO�8Y�ҥ����2��Iy寥�A�(R�HJ�Y��Ks��;\Y�X�wv��nT��w��vF7��̜U�v�Yk�i75�}�V�O�񷋽�n(f"�s"�����N[Y�U���*Hg7�fV�Ϥ�un��E��~X?6�e�~�
��;��rK�=:S�im�F��{Jf�ב.�)��.cj�>؎�Kf�}�����2-)4�sWQG���d�����=&��w��U�����m�Nj��zkQ��P����7�ٰ��H���V��,s�^��Qn���ʵ�c�n|x�Z�fM��6��g6ٯ�WU7����H��]Q���a�"r7�% �e��kԂ�FEa��E���w�Z���N#�VFڃv�.��3����,:�%�a��Kaw�}�$&�,�-8o�J�9ݙ��2��N��c�c9ƈ�s�/)�Fj7/�6W�X.�%E�y"�h%�d1H�f/,�o�!����<�~Y����ܶ ��.�W&p9-�R�P�)4۱��:s㣩����-�O� 0���Rb��`߇��*���{ఙ����OE�훱�8�l0���*��Q(n�߹f��-�tl�..�f�N���#M!���!��r˅,ˉ������)��nDHQ�sU0/৑:�z���~G���\4����烊;�1�4��R<L��}�;�X������^�+�M���R?��6�W��^'�\G^�R}?<�<]�fn�%*���T�AC�)1�_�d'��O�K1Iq���ʩ� �C�a���V^�k;�Ҩ�@;�d�����J%+9�����W�5HT~ޤl�Y��}���
u����RLqh%d�\��唣
���{\�����1��n�E|��$�h�`6[`�N�}��i���T��q�%���c�%�{�߳����)S
B��2��Zj����9�/�6������?�
���#���5Zj�8��PR��+V{�}6�ݟ�*� �È��y5^���d�Hۮ��e���y\�x�-:�Ӿ�Y�[7����f�D���r�W ��C����H�����2��2���_ewƗ�ۗ*�QxS��~o�]�M1�[�6�����]3����N��{H�$���6����`�Fy���B�%	��h� cl�,�8��!�V��H��f4�����~	����Ã��zh������zO���`=z���紗��x�W�b���d�W�*�,�"��V<S,}�]��ԶB�~��Q��[�O:��8���\K�����#nB�'m��
���P�3:N��#w��[N�v��/A�#�R���@�p39e�>k[7ԟB�?jB^�ǎ�=�͡$�S:���r�4ݵ�?��ߧ����{r��Ȫ~{@��D[;h�ك��)� \�����fS��@��[e��wA�.�e��č�M�O�`98��j_�m���$zȰ�I��Ě	�&���9��7���%�h�0s���Z�lL^�B2Ƭ��Y���fx��m��!�V�D�FG-L�O�ie�C1$��`Az�8����Ԭ��ˍNt�Q�uٜ6�;iRe���e�.h�J �08�>����D�^��a3{�������x����x~�{����,!c�kA���Y��HPmƺPosd|��$��≽Dr9������#��n�E�����Nf1!g%����st��{2���HOr�� R��*F7�������߿yw6]�iPQ��<��Et��k�ƇK*z�;�1��]�v����4�=�3�}�DoG�;dAz�z t����0Iz�v�L�����Jv� ,S�n�BZK/���}7'�^~}���u$V]���b9?��y<�lɐxpr���c)��Y������~[#��� X	�)aÞ�/��A���m�w��8��g�-���/$��Z5H \6�J���3M�C�X����q�}b���S��g���3P鍩���Q��'�'D	
o���oi�hԖ�"�@F����ҹ�w
�)��g�
������ U4V�
�&�w$Mo������P�'�B�����
O�HiѸ�B�W[��n���u-�	�P߽�}?*��>&���6�`w@L/�Z��k:d�J���4H�q�>/���ʋ�7,�!�'г��`��_��5i�{���r���k��i\sܟ��v��[8�FO7�evp��&%SZ�'��s7/:��=�ͼp��Hz���g=��fm���#d?MT�f5���Ј�laZx�*ƫ��f�S}�u2U�gƴC�,;-|x�SL0N^��]6�`���t}������=���\�ή�����Ф����� Tti���%(��J5��|������"�V=�$)�ᴻ���5�b%:��W�Sn?�!8醪������]R]"�I0��l���q%5Z���M*�/�%̀��U�����\f��*�������]�67�I��*��������2}��F�W����O�}?�"�S;f����w_M�.�	{�`J�vT��k,Ӝ=+s�������~,y6�42x�^'$M���/��n&��AB��X[�������� r\�ٔ��g�c:&�Vc��_Ju#�j�'�����1��P&��qǤJp��e�"s�]cC����r��A;s���igO7$��t�97f���h�ߪ����s�v�=T�{�,s2���bz�̵QG8M'ըf=9'x�I��KE�JR����^"�m.�PN㑓�m�l��@��y��vj�9�,�6@
$���5�M���jw��E1�X4#�9nw�ׅ��{����v٫�����U	}�?�7��+Y�䟩1�=�$�a� Ԡ]j�;�]��!�tj[�S����E��wa1Z`�8bcJ��B$h0}��� O��3+��2��:��L�M��x��a�n���pI
ru������4���E<�_P�b�����LO��1ގ����3x�eΡ?��OW\"� Hf) �_��"O-��T	�}>R6��9��zJ	|�L�ZW���W����g���J�N������b5h�L5�m{���U6S�K�]�Th�.�_/V�	e�KO��D:�AX���E�y��|��.�rW4d�D�v�`!Gv�7���T���ф�Ag;!J,���s��w*&VZۦ���s$�Qq`�ԍ�R$�)�
.�O��F��h#���;X`����h�t�4��O��K�.��`^��X��a  M7���0f�����n'T��d5P�3+x�����駌�]����S�3��P���/� ��~M�8P�'������N���n�kC���й�<�_ݖ�Y#A�E!�i��j憬�2m��f���ܧ7�p'T���Jpg�ٙ�ӐO<{����ƴ/���ȝ����u�&���c��"f8���N�M{�Д�Q����R����U���̒Qv^{)��;�$� �zsS�mka�����c�����ڎW�$|3�΋��D��W"�ib5�^_m��3ֻ�1DVy���S���)+{�K������Y�d�����z��o���?�!��|0O_��Oqqsk9W�W����d�M"ฎ�
��g@���vA�.΃О��\4Xu93�T-i7���t��!$>��������4L�}Ohz^.{�Y\������C I����0�T+�:�]���-�2�E�}�y�:�q���0�[Ȕɚ|�U�"Pe_jJ3���$�u*,���`ZJ�`��Z<���#��L]ߐ���Z]�S6*ǏB�����a�6�m��_���������-�vv"r�Ӧ!u�����W�`��̹޾�l9Ȉ%�0�[~w[�T���1�H�a���ui삅���V��3َG��d�8NE���Er�^��A+8H��{W	�?�;�VFӴA��M��:�(�(��u霾��<X���.�+JgV�|_����a�Ļ�+�+f������+-��!:����ܥE��G���%'U$�w4}���é�TA�9�L�4�$Ý�Oì�L����i����m��O��@)vz�����2f�f����kj�FF��Ǒh���)x��{�ud�zt��1�Gnߡ��J��z3�5�zz����5�VАL"Řw�̦Ϭ�{}^��}BP��fj��ȳSx���`�f������iR�c#�q����,?p�ԹÓ������Ѻo]�e>�'%M����M��E�\�dh7%���'���qLn�v~@j�r$^D��5����f~R�K��W���W����_����ʥ���'��}� ;�R�U	S�[V���Y��R�e�꫉"��E�t�{_�ԧ��1�J�
0ҟ0��|�u�8�T~b9���s�W�k�VI����7�<h��%~m�`�-��g�%�5-�:ut��#��0kj�"p����m,�R$�ʆ3$N���Q��RhEJ�O0����9�FW?�c��h���Ë�c���e]Ϧ8�=˘�^�#[&��c����e��Y �>�w���q<+	�=k��nw��DK1˛Q���+��ץ��~B�aa^��]����s9\�{;`ž�u6/�ы�f7y�"�B�N��;e�h]�3���G�1��ƻ����$%v�`e���
p!- g�hwrX�g]�E�q��0����x���s���b�'GK�N�K��r�d���E�z}�m*�Γ�[!;�3�����2gѴ�� ��X(��?O/��ؽ�i@���O`j��~��	�ŀ���*  4 �)[�qN�m�
�V���DĖ&���Ü�q����At�����ˠ�����`�z��� c��"`�A���8`��lQ/��0��/���i�^h'3���:���b��L��6'�Ar�U��"�����e\�y��v�.R��~dL�`��Ƭ�cMz��1e)��ò8�G�*�,��{ݸ-�����3���W�ƊP�5Ŵ�dH�uP��}�c�fz>�-�� ?OzU�� �T?1`0����Bu���|O�ݥ��j���3-�t8�E0i.�oX����E���HJ^��><�cR%3(SƢ��0���BHﬆ���o\a���}�[��q��Y�¸�ߢ�Y�.�'\G�q6�q�gO�����*��� ����i�v1��MU�`uo('c�5�Ak�@Yc���r��,�\Q��MM��������w�>�G^n��,��#���-"�¢����O��A#����3����j�^�%���i�-����J�pk�+���g�v�A�{�,5����b�$������z�����ރ\_��Iz⏉(�p���7,-dǔ��u�U��`��������`
� y���Y�T��Z�i�1���rb�x#�g�� ����n�r��O��qb꠯��dl@Ȯ:
-漸��o������U�p�ɢ�K��a奙�F6m�hoXbP��0˞��T-"�ȩ�����>��x@�e0��Q<[,��f����>�Ƚs+F�0����n���(*����'��]f�/tjs��`(�$"�RF���N�b�o!rt�{h�Hw_��
K������3�O�n$m����/�[��<y �v��Y@��+��:��E[2c�W�0i�����K��*.�7>Y�ad:�_E��?�i�!Ʀ��������
& ꢐ��=�٭N�� C
@,�>'��#�ELO�gwZ��(�f�T�e�>@?�w�~�Y�MY<ІH@����O~��찔a�jYRij�K?���L���ccU���|��Z|��w��#�ށl5��f�8�7���7�8	c�)̓Qp��.`vO2k|�vs�{�����Ο�s�v��5Bl&͡�I�\�UI�*\�!2���S�#԰�Gabw�V�K���G0۵I����x���/_�����ɋ��c�?BR�d��%�1�t���Ѻz�т+|n���}A.�"ׂ�� !F�7ӫΚd����>��=n6�&`%�=,�4��p��y��	l3Ad��Gh@yh��9,�sY&9w8/�E�P���j�XSo)�3�3�(f�F_�kH�R(C��A��`��2o+5Ω� ��#}4�ۨ���+���x�Q���������k`<E����^�T��(0^Yo�
)�W�T�Ø�P@�r�� �~�&��E7ӳ@�4���-�t�cQD`�X�/%��W��k����e�e	�/�Ҩ����l�se�Q�0d���d�
tSk�|��v���,�j�>2*VE��B�#�T[!���n`d�3&���lr�Q�и>�E߲\�M#A5J����=ȉI-�U�v��#��5hOU��X\�;����3�����`��$���'���<X��Ҿ�a�Mt��4ӈ��{�jLe����-^�9�\��k�w��5���I%�UlE��1��I���8o>�)X�+�}�|Xt!TI[�Yi԰��l}��K@�����N�m�\q�j#3�>Ʈ��UE�(�oͽ��x/���*4$�*��!kQO�E���<Ѧ4�����K)ӦK�v����]�1��}fT���Y�&���%�J�B�&����4��4Δ
w�{�+�_J���*di?�9��!�V +�vV��3�=��S�p�Ե�,���������� B| �7>h�+�)$!�f�\�9(d����s(M�Ο��1䬕���a���%�ic����K�KPH���!S&׫=nS+y%�5�� ��	���j�i���h�{t]�������B*�۬�{o%��Z��-���4y{�C���H��­�?�����g��5�J�Q�X~�EZ�������!�˒ 7��%�X���hs��ϗ��x,C��O�Ä���^����*�WH?�,
E��`��_�a�@��@ش��5�!$`���Df�����	2~���+R��ӆ�O�KxS��D���Ns�z���ۆV׹���B�LII�X3��o�o�^�lAY\�;/A�t4�ofG�[0O��]n�]��{�E��D��H��xauV2����}H�K�z�~�j�䭝�o����������!υKS��q��[�M�̛Q_�����O�@�Ӏ���EQ*ho�8`���=R�<f`Sv)��E>O_%�x]�V ����Xx xߎGW�UX6;���;z)��#��rY�`��'DG�c]ڙ%��
F��c�s˓�,V*��,��k���m0��V�4�]K7��l�����avV`�${�}0�%-��E��� �h�>�D��8��� dQ�	>���Z2�̝����(˯O:�5�P5���@~y􀊝�Z췯M1��%'�Kٽ'~+<��/��:�@�&��qpn�ivs'��?>/lxO�ͱ���Q� ��K֑:lS��rq���f�1͸�o�A��x���T���O+(�|P�E����LX5�|��3�h��k�;�1񭍜�)߰&C��h����!JЃ�!=����J�p1��7��E��|,� F���>4C_����7S��i!��.���.xw��N��&��S�,�t0Խ�� ?�_:qň�g�������� N��d�@
���[���G��ݫ�3�D��62_'��/E<�1{�������͍�E�B3�WĄ�_��P%�<<�!%.��FXZ��:c�j9����\�z�SX�)����-q�sM�L���WcpQ�?La��g��w�؈�Z4�l��ў���:��bu�bT�M�V����<f�e�d*=5��,g�z�5�M;�'~:.;�E����FqB��p���je��j��+S�.���@��Cpm,���ٱ&��L<r[<l �g�4�\���O;?73�%������Ak6B�͟=dӿ`��nȹ%t���C�C&����k�z	Ajɠ�1Z]��>��c�A
δ���MϲOp��1O�3�R��y7(�e��_K�j@b�귑�|�����T�^�;��OcN�&�Zn�2�mp��-�k(���Z��ah\g�� \�.J9����;��
b��k@� /M�"�	��?�/#_��nY>5�u����x�%,% �?jt����]D:�Lη}��o�-�\��q2�m������o6{3�9�N�|�7��K#z�� ��a*���t��πHF��n�j��d�\�e+�����hj>���v��6O�I|e3(������v��Il���� �I!IDJ_h�͵ĸ�G���%��WSkog.��g ��o����<�r��lk����/�d���#\�I�F\�cd��m� �l�yKժ���y���~��'S��&D;�=I�����n�b�cuc���0�ZK�<���w��l����`m��͓����&S���cj/�n^�{��O��98��Q2Nk���?(�_�tf}�=�|j&� ��Ap�J��tO3���������uL��;��O+ʇ���sm*
I݀�J�W���A��~ʖ7O�\E��.!'��|��/o񠾁O��
k����x���[K٪M�I��|hwfo��# ��T*�ǣ��ϸLW��x3��s^����a_K��b��k�L�Q����!5@}�r���N�Mt�7�?&����nU��c+Y�#7 ��t�qIxq
�j����V�g�k,��n�bW�y\�S�f��C˫@��~�#Gǥd����IbF.���0��W��T�I�'Pc���6ĺF�=ˡo=�� A��	�P�ø�P�ù�H}���7
�F���7Nc��BQ�?Ho�+��k�Fa�);�xK~!����[�T��$&�#�WL��r`��~�Q��/��r60c�����m�-1ҵ�B7T��Ƀ�8���1�l�ܦ�7.CI�C=��0-�qy*�UO�vr��KҨ���M\z�݇`�kr1T ,��eۑ��m���}2f%��WR#㱲I[$��w���'T��F���a�;����Vh��&���v��11�2����}D��kp5C�p����-+�����l�NR�Z�F��y�� ��}~xce˳�8
s�t��~��1�K�l�dJ�96�7��~�����|�����4��	�� ����^%����ĕ��D#�!� ��ǟ$�����$*K�+ч}X�T0��hY$��7�<��y�?^�ρ���a�".�9!
nK��Β"Y)�;{ǇC�P<؎k���h�1=�=n}�ۿ���F�Қ,�M�R�v)-0y�<���;�&X\��(XU0�� �F։��l@�CA�a+U-�7����6�ϣ�]���X�lk��q�f�
ܻnS6�?v�J�&6�����CIB�0��XG1
��,�@�s�n��ٷ��	��]g)]��O�b�cb]r�#EB1�!�ύgֆ3�[E0�+8��V$�	0
��sl{���hbY�o�� �Ѐz��v�A:����G��n$ ]�2��&��a^ə:�b���YY���?��ƋE�Q1G5�f�<�E6h �4#��;��0�i�&���\Y�Qͤ�~��e��S����	ג��^��d�9��D�M2$��m}�O�*�ϵ8/Y�������w�T��J[������Ȝ�O�q�ϡL!�7)C|�
�w�*�ihSڥ��J�+��ei0Mjs����W�=���ҍж izYd)��f&��E޵��3
_�#[���8�v{,?���|M���m���}�����Q���&Vl�\�p�>��1����'\ID�����7����	���� W37�������4�XIԠ��-� k����i��X]���@\o�H-���e�Wkr��d`�jXT��4?u�We0�;b�-��B��^�-�?@���J�)$AvCVUd B3�}]$s*��VH�nB.��I*�E/uY-�;���L:@�{� k�kFe���AǐG4���5k�W���m����T���m�ȼE�?����);/�ɀ�3�}{��}�N�b��x�z3����!���P$ɂ�N�ܖ&l��%9.�N�r�ٛ��f��F8��5�d1�\/DR=SBk�;�?���]|��S�9�`B>��e��Z��~ھ�C�%��`#���d�������dj�ס��;��5h~��Wde�=H����`1s�"O�j�ש
����{�0j��D�j�o�|��Px��1�[��e/�o��^���f2���x������6�ul[F��&��v�2��O�aP�ّ��c�
6��Nޙ�пmV�o���:}$GƿW�9DF������ٍtP��Ӌ�JE�f��,��~������ ��Nf�6�������#y�VQ����P��F"��ֲ`7���(0�-{]��_g����v�Ç0�%d���UM�Hc�����Wa
bý����W@L���m��w^�$Q��Q����e�1�*7�I�?׮�f)���zh-�J+g�d=.�l��G��#��F3�0�E��<�P[�jT$,Z)�0)������u����e7���jg��Zbޔ�F�r�d�ʮX������7�u��4�j)��X�l�
��qi�&`�<�c��}e�����Q荐��ȇ"^~�NLr����Q��{'wE���f��)�͔#�b��9�V~��@S�*��GP��#�2�K���p����b��xH��	��uԽ��=��n���?��5�`1�QS��;�}a�[�T^)�g�y�ʰ�L�(Y��XgeK�{aE�}�σ�6K��P?��Mx|-X��X��|7�>���g~��ó?M^%�3﫻;Cm��RɮC_~�E9�8 N� �/�T��R��W$i��s�
F�`7��ZsX�1��sR���cԐ��mf��.����%w^e7I��.��7݈y�v�`�F<Hi��v�}U�����wf
eZ���(�~l���̡�=�h��xCHa�Y�vu���vӶ���SOa�~z���= 6��@���W���δ�
���_ԯF���\�$�E5�8�G�vρ�9a�OGp������u��Y��Q�D��#����8If)�P��`���>p%p7G�T���y���YԕE<�m���6�s߀[�L���!� �Г���7֙�nm�l-H�5Ч�r;�)+��?FG_�|���R��l�iv�$�[���=Z�p�'AGa*ص���Z�LO��#���w��(uë�Z��7I����������`�c kE%ࡋ�2}|��oU��5\F\6>1lq��bi�:أ�{ϧ	=��&[S/p���&a��zجq����i��'�6��0�r��.ܮ���>�k����sīܻ�:3���q2<|A_���~&<4���ءKy
�P��=?����
zy��D#>��kudx�}�34H�"9u9�<6Ip�@�OJ��+�.�xk��b����㚹i���|cS����f	��7��F�__����ʦǏQ���׎�^���Ϳ�Y���Vc�Ѵl���Z���=�γ�q���_j�EG�Tl���dU�ɑl3�3�>ҍ�d�s>��f�n��17M�ВEo^ 2�ƣ����/~���d+�.�4H�v��98f:�([v�\b��B���ͪ�yB�Qm�y�=�c���v b%�w�����\��>C/SiJi� O �ɋ�3�UV����"����]�"���e��n�w#�����W�����C�������:R�7-��K������
�@:��a�&z��}�3��꿁s��;�;8,:�����?Z�?%E8'e��y Z�kN�f#�������C�9:�J.e�\�SW.��
����C�KYV��9�ϱ��S4�{}"4�3��� �G�@��ҝ�����:1��aj�u�+^Bc�d���lI)`1!�8P|~1*~�-���P���7G��t�~X�<r�%IE��i�J<����~�k/��H7M��"�'`9����c��P�s�%��Ԛ�CJ���M�}�1Lk�]�b�Iljy�-� 2�p�p�w1�;��XF���Rٌ����C3�DT�!@�XU�ld���g�pF*��.����n��U�@��m�c�~��|0r�J�GV��c��&_]���n5�׈�c�x�Q��!!ecE3��ĸ*�i��$n��N��q(|8�����׉��	�,�C?]夳��/c:�zڊ��J�P��.a6��쭎cCI��{r���&�E/�x ;uw[��4��8�K�4�[���c�,&�eG#�&��yD(L8��j����kMHպ��h=`������H�p���SW�S4���y8I�_�e�^D���5S�!��JRlQ1
�� �Y��z<�ԙ�(�'3%����؆�B��B��h�zcѣg�Ψ�7~�����<��/+��*�����T>��O�UqţK��*�s��Y^i�=��V�T���&����mBQ���6�K�s��fW5#T&\��dKˮ�5�D.�jk��`9�؀�ľq0j��#DL9iQ�*/[�Z*�᝟�C�5[1����+�邔N�Uw�\Jy_k��R��<~�?lj�*��_&��w%�u�ݤ��%��"Ú�ȡI~��~��]ZA���l�Ӛk,���K[��͉���׼��@�K!��#�3�Y��U	�1�Ә���j�ר��(���d<�w���}��$��C}{���0�]�
���� ����0�Q0�`��u<����1�d���yi.Q.~�mT谼-m����F����("!\�l�؋����a�;����.���ǉʇ��g�� �9e�,�����^��k�m�H���楶��	}y4(4�Jk��3�B�? ʸ(rh�:�Y��?��-��Ġ�[:�:�t�h�?�$�V�v�u��=��Өt|AAp��wph��ʪ���ޭ^�S��;�_s҄��b}� |C��06ѯ]=�U�8K�ʠF붳_��9N9W��i��U&��~�iJp�څ���&���*m�X(�:kAI���AC{)�t���6Y�&9����.z3w%�ȇ2dv?V����2w*�HP���B��řH6LV�˵�G��x���e�=�?���!�V�Y}��5Z��K�R�4����
>*�����G�:�؏�ʮ:�4#W�81��L�/��n��k��^m�] �ׄ��q�37��B�q�q[�su���.���l5�ٿɑ�E��qsV�w/O6�\mawH�˜�h��zr�L��f�N�lI1��d�I Ȑ]�<�L!z�=��<�Mf�S�RŔ۔�m'��4n�P.��a �Ŕ�zƈ���D�&^y_���������#zW��@���1���'�Y���5�qft0$�B��V˄�\~B�Q�Cu�)Iz�����?���t�yM��KՆz��|B�w>�~����'ʭ����_�j�F�~��'��T��$#�����L�c`3��q�K��e3�)"�S�1+Mg��؋f����O��[s���R�:�N�㝩f9�@z^���H̈W(�u��ړ����U���x�_]�Ȭ�E�@\��V�6�D]�Ie����!��P��G�)ܡ���O�`�o�34�$]춳�H2_.����Z�<��G��#I��.�aywڰ���E}���Pj��/fI��QIP�� ��ִ^�qA�MZ\��)����:�/�c�r���z��fK�x͘ m䴶mw�]��ωr+j��Wyq-��G��C���>���h[p�u�F�ń��n��	�@ ��H7�RWeŹ�E������E�!��3�f( �'WW�<Ų��l0c ��^_¥7�g2p#�twA[���Jb�C �*�U���a�o�-�rR��j�Q&���+�L����'e<,�<�#7����u@���=\o��4�Vws��e�&X�r7��M�s�մV	Ў#��Ԁ,�=� Ϧ� ��07����ҿFa|������O��DB��Cr��b�.�b�����|���-�׺��r�0N׫A�>��IL�\��5D	�h�O��V���J���(�h��쓆�j��	�B}Ꭽ!t�����tAkC���OU�!1ߖm��<�ǯ�WL1�1��DPi���^�U����}g��;/u��ewC��,3_�кR�Ju�=	�	ϿT�����ԥ:N)N�m�	M �: F������^�Z*,�������N�'aC��,.Vu�b���z�t;!k�!ѕ�zQߺΠ.^�_����b���!-���+!�q��VÇk�ޓn��z��:�l����<�>��~��]\��| �����O"� ¨���h[�Т��%�l���zlЩe���q���g,��C�[[���4���G�܍QE���Y�u��%,�7��1G�y�5��BK��mJ<! c� ,;�0�Z*{.���>�Nn�R�Dî�[�v�NdV9��|Ik��ț�/-:F�qV�`�c�5����K*��F�����7�ob3�P��r ���@�M�a״
�������\��:Q�F}@�L�V%�{
p}���,�H��/�e����ɵi���F�ߑ<� eZy�0��\�Ҡ�0fi���i�����<�=�d��-�W��u�����<#���H�O�\+�p�t;�jp�"A4�x\��#��%f&�H�Cm9>�mB_�f�q*j�)��̩�Dr0�	���t��Tg������2�z�H���t}-5��d��t��1-I����S�?A�d1q�H����3�����C�AA4ORE!��Q+'-U�d��҆����S�"i���{W��,,�5g^/����i��r�����A��y��_���@A_�My3$F��.3g�M�}5�.2*t�q��5���	۱z�$��gp���Ri�+S�G��^җ1Nǭ�5W�a�g��M�adbC�bz����t�����U���ŝ�����~%�FA��߫ c�C+�A$��!������F��,�[��F��	����ĕ�ߧ��u����{��==��Ir��ˉ�L6��N�W�ꝉi�Y|��k2��V�M1�VZ?�k,���+�rC���K�=XAE�b!�(b2gJ�e�	��ï ���A�'3�9#��	oxh�ƙ"h>/W�D)'���6���0M��o�[�8�r�^Jm"(���'����?�����hԆl5��J�1�2�c�^�b&Mg������ۆ�v�Wo^y�i�/���?��I
�B��W���_V�_����u�d���Jf����Tg����o"�ι}��8���n�?\�Y�O��+��;�Y��[�˶�?�ｅ㿘;��@�Ur�.� ���>�|�Və��%�NF���F��0�,e���S�Z��\>�`-b�S�g�
��gp�ǹ�Y���в�wD��5Y�0OTr�)�=�F��J3r����(u���:�gԿMgנb�*A՛���˽͒����w l���S���Y�yg�H�m���Ã�vB/Z&�&��Z	�K@�Z"sY�m��'y������I]�P�ʳ�O<E�Es?�>�ɋW��Xw�����0僊�=q"z���eQ�NV���g�ך5P�ډhԘIT�=�L�X*鷞g�l�� ��H���������#��={�?�jA��B�:{U�](v��<��U{*T�Ɋ̋�Q�a3&Ӷ_H��K��)���~;�����G�X2?D_�65�<G��9^��� O�g��x����ze$�l�a�zN��3	gc'��[%#�2,F̥�����V��X�8�4Z�m��������0�S/��#t��J*��A6��c9k��jNK�(��f-ju�ѻ�فl��5o{HR
d��_eAYS2أ2�'����B�����l Cc��pEzM"�R3��_"������4����}�-ё�DIi���Y�� K#e��U�\*�|�U��@�g����]`�����a�g-� ��U��w��D,�&|"��~��i���^�I�͸�D�:�a=}�b#�ƺڙ�0tU��L����`���,
�O/s �|�Y�W�'$����0����ܩ=�#��=�w�2A�i~rׇ~��.��Oi+_�Ng���+Տt��\��ȹ#��p�#���}����	�a��@���dh}�
b�g����uG�3��'`��<��`�6��-ZC@��a��Z����M�ꍎ��l�S,⽌�0Y�}	Ƈ7��	���a�Nw���1�*f~|��P�x_��(�¤-��M'p�U�f��f�^8��P��
��P�k��-x���t���ݭ,g����b��_��P��?�O�{��F��w��x 4����+O�3<O�z׾ԁc]8v�_<��ys��Q$L鱽�ũzN����"�iV�9�6p*���>���G��F�)��8���U��jn�>�gT�۴(�Y<�B�i��*Esb�e����r�QFT`$�ɋdd��:0B��Cآ:�K���!w/�!4P�
MԊ?4�'j<�LnEA�X�_>��>?G�7�1
�
zQ��ޏ�aF���~��-}���GOV�:�~�y}l�n-F�!����ΞHI
%���%��)�]���+]Aѩ8�MV�������a�a�>�b��E�}V�h �/8�F��I�2E>KF������~�aF��m�+�d�n�NT㝪/�,S�'�� "y�`H��9dEH����7�u��/
����;�")z���P��s �hL0Gz���q�䛿¼[��'��/�W vޞOF�˩Ty�jU/⠝5�����I�,���wmj����Z�rF9w_�� Skb��xc�x���Q5�� {���5V^������xvb���K)�˜��������*k�j�n4�}��ᰛD����Nx�W���o�c��NS�Q?�e�N������L�Σ��G��K�l\4
�ǖiO����]����:��:��Sa8�@��jP�O����Jd� ƪ�:�K���FM��\Tg*m�pn�9޶:~�[X(Yv���d�؀���Bp輷y]� ��T�H!X�U�����z��9Nfn�n+�Y���(Ro�L ~�am�G�2Sa
4��sm��~�'��K|������{ʂ��)�L�T��v��ҿ}��}�%�I\�<�3&!Tx6��V<��|������o&��J�WD��;�2��<3���zC��wP�q�r���M4��`�jK�CY�����m�I�r�E��}����ҬJHGTD?@-rK�t2 >7eY��|���������M�p$����VW0@6(�$���� ӕ��w~dyQ�������aӊ̂���Y�|��8]u,]��qB���G|F�ǻGk
����f��U�vҵ�������X�絒g��>?��1U sş�*�^��0h�2J{i�t��u��bA%g�Q���s���3�����g�좹xgA \���^i�4���#�D�ed�z���
��[�*Q�N�����h���X�^����Ĳ�bH��C�F�D0߇b/�1"A�G5�|mjmN��v�_�$շ�/@�]G�yv��E%�A4-�jz)䓍G���=;��w-���y(�pg�G����z(��f��	O�v9�h�z�I�Vt��[Hr ��p���'~>1 ���W*������,yv�:�t�"�X�N}���g�͌�x@Gڳ۷�  ��rw����"��d�Mm����p�Γ�}�T�E��@��#H-^��e'"�ޖ��2yO�<ԩ��o;`��P���݇���I��W��޲[��L={!�	�ύ��!ҷ�,v�Ov�+i� T
�4�-R��7�j�X�\�C1�;�5��Q\2H�un��b�M� ��}qr��D?'OQK/r��{�#g��hR�k�7�{Rg����Ik����u�p���e�n�Pf�a8�	&���:�IP�{��:�lCy��t����Z}�C�2��m���MZ���TJSL�O����1a���!�}�m}h���^u���"��,���;��4Xi8�htن��2�F���F.ϱ+v��m`�v��ģws�8�J�҆Ic����v�H��@=yH���#��k��;,~�7G��T�rz�������6}s���G��%����k(�"�J��}�Oh�|�Q���O�tJ�_��}�e�lɭ�=�v�O!S����XpDэϗj�?����۶���SY�F�;���:�����ר{}GsAO�T��g>|���V�ઞt ���a=����	��_����2 ��Uj����c��OeCy��u���m?%�؜@��E����9�T�n���<���FV��<�Ջ��,�_���4�
��Ð����t��Ғ���;ic�jUPI�u�qO�x� �eŌ1�(��|Oε�D
[e/������'(�I�EO�z�p`�/��d	Y��wJ��b-_;��?�A��]��cz��{Eot�FX�k0*1;�yTƜ֠�l�ͽH�/���S�4N����N�oQk'�$�#��)z����|�!�fPsR�H�:DM�����Y8�{d��x�k��Z~̻�zc|<�PC ��mTvs�p�������lp�ف�k��H��R �p��Z��h5�J���Ђ|�)��~Y�F�z���kd��)���]R��[����T�P���O�Fr� �O�gS~�/V `Ԓ�����e6)NZ�}� �:>�ˁOHa����#��%���9X�D��znO;��f~�-�ڑޤ�T��y�:�~6�1�Qi�3�05���H.�"�;�4���½�B��Ы�x4Yr���Sg[�X��X��[?����h�)�G%����agz�; ���Ώueʀ��;!Mq�����kJ�'����r���ϲ�Rt'.� #T�����LT'����E8(�PztX�B�����l����rڹ�/ٝ�v��K��B82��X��'����Dklj�S��znZ䓍8`P-��%�o��r�.�����V�ǊH���ۏ�M�q������F�fd�nV:�!�B�ɟ����r�QC#~r?K����W����>O�`�0�s�T큋%�����~�o���o��$%�۴�����ܣ4��+�L{+2���|x0���=�/�PT�ryX��wGM-R�º�}7�^�I����U|�  ��d�z�1�/���ۑc�V��w�<KR���V�+�`#���p���3��T�7��a�c�"���W�M�	l�����4x���7��� 9�:�^���,5�.�9˛R���f��e�	�l�Ha>�Ś����N���BR�2�ͽߣl��t�\ox*�\�-;-ف���jc����K��&�|�]|�kdC�r�ə�M��BDĖ�l]���o
��~����!b߸�z�>U�x�����4$=�f`~�Q��ߏ�j�=ܣx��M��D�̘�u���	���/5��fQC���4�JA[Q�=) &�&g�"��cً"�s=u�o�n���J�����r�y�s��L�=IX~���~��[b����7gP��B��v=ΟDl~z}VIV�����-��C`h=��O�N$�L�IQ�ѷDMDU�>�	س$��n4��M��/�l65JP�� �N4s�m���v�����_D6�x���<��������w�Y�pEKOb�+���r�\NSmM}\����,�w�%�.U3����u;>pd��ʽ>\�7E@|��p�|�Y�"�]C�#��Z�䞩��ѡ��v@�/����Q�����͊�Ic��w�r�� ��NI�T�Y��\�o�]��/�G$zO����:�"+�>����F�*��vl+oF�����c~��a �͖$�Q���P69`Cr��g􋣐s�̀Z�Ǖ=��5[��L�jT��"}
�@�V��M%�"��(�@ռĖ,�����sB��a���V����쳇c}�}����a4�@h<L��V�����M���qv\��v���8�?�ٺ��ג�q�PF?د���ؔ9W��B�]��m#��b la���$�C�!��]���C�q���5�2��T��g�k[�[�����?ꭒrX�Q�h�)Vc�w#��KFz��ۆ�UFJE�Թ���R	�����+�_8�P$�� s���2��j�S��dl�5?�e$k��I�WG�E�]��.8����co^ehT��i�U����E*M�'a�FK��k־X��m��W��&�2p�!BԽx{0u�t�ZUJw��?GF_&�Ӈ��]���*<9B!8����1���`�Ǒ�T�0���<����6��
��^�/������W������[s��N}CƑ��AYl`�d-�-�꫓��|��b�@�Ƹmw�����	���cm�R2ռ��BM;B����vl�MK�Cl�l��t(f$NN�n��~y���� ������p4�L����[PG��G���@�;����dU(<���R��v$!qb��z{U�iD}�+�zz��@8��X����Xݼo��&��·����OmV����E.���-�coǈw�4��m�婚���)�s��CMQ5�O7az#�����~M>�]c}W���Qߝ%�7���#�W��>U��g@�5�>�U��.1 52�6I�չ��:ʶ�*����M��e�am���y6�Da�34���+.{N�-��:�z�]�����٦-�v_S�${���U����Ypm8�Wor4.�����);��+l��e�l�ֆ����gѪG��7���L*y�mپeK �~ v��tX@��cS9j�W��}�&�>��:D�Ɛ���C��?�*)��M�����LI#�H�	�|�;P.��?���)w�ߦ����Rd��q��d�!�W��4����&|�;7I�,��rn.��W�G�����:WGC�佁Ԓ��5���2$0@T4�B�zG�{�hL0�9ӯx�k�I�5�k����1�$%�%������$��,d	��?�5�,���!!�������W���x�mK�ަBM�� OG����ԉ���:0YM\���B�/?���P��8�V\�=�h��Q=xЭ���^u����}`�M��A�F6n?��/6ଡ଼���NՓ�QΈ�Z����g$S�Q����ͦ[
�*Fd9�Y]�;���_M0hhr��TmѠ���t���� ]�EwF��䯥
)"��.�%���M�0�m%*�j��7	-�]=�5\�Q�y����l_�*����w��bAa#��U��:L%��lfǈX}�4[M�9���P|,�;K�B��v��7�`5�"��V�%�ӡPn�sۜ����~o41��Ҏ=7Bs�ͮK>�ک���t&�|yI�vCd�g�#;���?g���D��7� �o +<��(��R�Ή�} �������'#�p�gZM��R��f��PH�H��&خ�fX"�0��]��$T��SέD�2����!v������xN��p�Bq�� �IN���;ֻ����c�m_Y���ԠH�S%T��@ZԊ���f�.�-�!����4��dFJrкاi�w[O�����Φm�qn,qB���Q�3,:���z�db��S�wq�3��T:.��`ҔãØwD�I�N�����dv2�m�����~��CJ�UrnZ$k��d
�����c9M<_Q��1�cO�ґ���s� �V�ħ�yZ&�i��[��m_��l�����s%����V��;����<�@�H���D���8i�0?�;�+�!:P���n�h�j
U0���cb���l�I���cj�<ϵ�јxė䝢�ylMEެ�/�b��JDA���x���Z��J2�zՕ?(�f�V��@Lr|��h:Em�8�����Ҏ�F�++�W�x��K��Lft��-�X�R(9�A�V7J�(5���T� �푫��|Ϳ��d&�IP�11tî��aȼs��:)�k��v�&"���[8� 'r�9&���k0�^"�пT��^�2��ȵU���9R昗��4�ǭ<��J�]��m�d�ϩ_���V�6�q����9`���0W��,t�Th�ܟ���2�mAA�_~�P71G^���D7ԥ�N��nDMw���{�b�[�yq���M&���/��d���ɽ��Q�M��Rw�Ą�R��p���\h���g���˜.���JKc�+!�^���Ԃ���d@���o�P(uwJ�#�ɇ	[����7͏���� 5)�H+-m}�'Q�6.������3PI�G�%?P���U�N��75+�L
���疗Mg���Z��`Ñ!^ ^�N�(�E�=pVh�č��6�ĵ)������] ����S�1�D���$T��Y��7c_�����5)UGS�%;<�"��&"�mW��Gz4B5����K�h���1��s��;��U�<V��݁^��P� �I��*^j�yj�!���{y,P����J������;����Ka��`qJS�Qa.�U*��oQ�"�,1�����m\)��`iz��\�,�����,���k�rJ�\����������y���!������6G���D��T�c����78^E[x�<����)wkR>��K+w��(jn�T�R�ȁ]x�]Y2�+Q�b�>U11��	q���	�5+B���Txs����9S����.��-oh̓-_P��B6�Ԁ�\���p����en�,z�x�!�2# ����$%Y��-�ba.��h�-jҏЍ�1�5���ߡ�%��&u��`�j��X<
���(�=6d<@9�㨛�*]�Z����el+H�Ӿlc��N��}�����I~����`���W�*g����ZU���3},#ݮ��/�V􋕒���*s� VfY��G>z��kH�����C�
kX�x(Q6�0�\x)"jL�*L# �OTM��Ws+�b�(3r2)�y�Ȩ~�t"���[Y��$����ap�4���Dq�+�)r�L��'���rBp�u�H��c��ZA���g[\ʫ ���K�-�S﷌�ь���n��ʻa�������x�$7��9|n�4f���yس��P�����������f��=92:��j�^C�[��F*P���3Q�P��f �
Ƃ�t|f)&s�:<���)4��'VM�1��Oe(!�~0Vh�~5o�ت,�=�Z��,�����ޕ΁�����iXUޚ�)�E[ A4i�60oT�Z���x�+�ͱ��cp��Nl�s�H�E�K�ru��$��p]��wC��B���l�x +��*o&�T�b}6�R�"�5Dg��`�dmZ�L.^:O`��Wp����n�l:"��(���y}i�oy��y;�Pp�-���@]�|U���aU��h��B�	w[i?e-t�)	�y����F�l��-�|�D�P"�ge�f$a�;Xh��fY>��$�S��J� \���vY�W���ᣃ�J�F\	)�����Ĺ��"�4����I���#��!��[��$wiPF>�{
�~����J3�����/��j�&{��3-1���2 T0s�.1��]�}�����4�O���`�W�¼�l��t�m��-��̸^�*!\��F�O��Ի+
�Y{�y���	�5�����?����iM�+,c������U��M)Z�4Bt�=���%�΋��
VL�!���_޸�!l�# �s���;&5��K�		u�nBH4�����y�-�[�9m�8X%	�[����\�O���c�cNꍦϧ��Ba�ӽ[d���E	���&��GY��]�v�-Dc@+�w�DE�SZ�9s�r���KW�o�牢Ti�k��W���K����J��s7�o�\��sւ.�[�H�&c�D�'�	��g��8�	A�����T��_F��|?"���Jd�8�K>��=uofF�TGȮ�쩄:sK仈�=%�it1�CJ����VW��nǶe���9�"N	s�hJ�:��sQūpC�E�a-���=Ts��t�D�p�NYj<#���T<��|6ЎT�Lw4�+��Ee@T��9{�P9OSb���\��,aWmk��I�uam`7R^5����,�]���n=�G�E�����|oʮ,����_pG��:�<ht���z|�>�rT� ��X������OX�%����I,$`Zڭi#������EN����n�����!rBS]�$Six����3C8|�[	n)&��"BY���+��!�ɒĳ(��b�$=��2B��Y�B+۶��1P앭�0a�k��6Ǹa�!��q�����2=���o)h	{�#���mI���<�%��MH����f���ɗ��q��N0�{l��d���t�O1�u���b��c����O�0v������o���֗<���^��M�-u��!�t0%�3�xE�u� ��@Cwiwv�����'Sf�]-��oy���ł7�|Z�ƶ�����%����]�/W���G����}=�h��-a�A�-��xm&�
�8�Hq������q?g8�"���
�0=���-��\0
��Ev�kL"V�i6��P�;b�;v��ၠ�"�͐{��5Hv�H�̗\z�׬ϐ@�?�)�u�[! ���)�� � ��;^G�p�h�#߯���� ����\x�����/���T�؜�]�~��w�p��s�[7@kFj��x/ �|�}�������Τ�M2�Ʌ�+����_C��2�rFpW;P�sxI[��RƄ?|z�"(�d^)4ǝF�	-���`��Ǯ?�,�:��ta7�z�̪p3��a�!_��ӹ�Y@�#�6r�x�vo4�lڎ=i��Q�+B���V\N "={<2C���p ��)��1⦤ۨ`�-�q]������q�3A�	E�+��;�����f��/wk��	�k�;L�=��gr~м�=R���񕔧3aDF�2M࢏���}��7�lR��{%8�$�.�Cf��
���l!�r�z>We�wյ8�I_���K��ʪ�����ٗT�N���(۲*UEl>�ƫu��SQȔ��{�?Ȇ�<Ư��ի��+��!��V]Q<�k4=�SJ��'�����.Uϣ�1��]x��3���L��|�������F�Rz�)��r�����IJ���8?Y�^.���,��?�@N��z���8X8�T�3l��GБ���f���]#SP��e(E���1���Ս��t��J�#��P"��\�r_��4g�ZOE�s�©�9���-�J븬
���#zA��r�Y�׮lR3�X�0b��m�m�x��r�⥿�*[�R�ԯť��h���O�D��A���e��8ZG��<(i�u_[?p�E��h݉�d�]�ߐ��7@�û�� ��e�v�f��y���wN��i��d�4@;٢��!b,�E#�y�5x��DB=
�!M�/���f�;(U�sD�O�iՈ/��Q˧D�0ٰ�ח����-A[N��g�c��HRF�*홴XɋsE���m��Y��2c�+��^y�`��7��[���i踴����Ѿ����>-8f�ɼl(����	9�m��J X������TƋJ`��X�g��p@��װ vʦp�<�M�1�gxѰ�̧� �9��� �l!��Qv�i�ش�d�i~�韋9�7����4259����j0�q��� �P-������[5O���3큃�U��M�u����V"L�E4�Nۙ#�NGoy�y�;ۄ�-k	�Q�rnh��S�A��g��*t:b.������Zi䓞J<���;?r=w	��q�F�cu�|��P�:�е��r�S�>a5!-�Q�[��H�;#rL0ʁ:��-�z�!�}[Xń�߈ʆ�O�眵������%��k��6g�?���;�؞�jr��Ru5�?����c+���n:�[l�!4�砗��@��A�o�1�k��-	Q]
 ��H�����	�[py7%nƃ	{|!���wj�cJ^���>sgz���p7Ԃ�+���B��TgH7���6�3P���ؽ|�|t����%G�8W1�e����/���!�1{��Y�m(&r��6����Cg��u�k�걕��G�su�-�Y�pw{
<t+,��3/��$&��ݘ��}���>f�� Ŭ9�H����w{P�]��W��d>5Pybˡ�p���*#�����m�J�h�搂G��4s�V�x��E���gw���3{)[���OܕƄ���U1�����L�����$aP;�h�:~�D�=F'���1��*bY
��B����	 	n�	�>�S�z���1r݀����,���j���
�����@߸�R	m����������ÛQ��[�Mf����+I����_N�����������I�#;n�5���~ǯ���d�V ���!b���L`��K�L;p�*���U]�9c�0�{Los��8X=�Kl�
L�~�o{ɂs����8?P�q�ͨ��s��|� 0#"�c�����l����|RQ��}���YW�ͺ�2�0�ͽ����ʪLF��g�7��;�'���ۨ��,�b������=/�"��/��k�I�g7��Qà��e���`;T��oe���\�E8�?�8z��?��M�z�l�/%��A�Ql;%�'�u��� �e5�&��{C��%Mi��$�Й�q�|��m_�=nk�\�J9�D�E$�݃(+$����$�@�w�-%%�p̌�x�[/�Z�r�t����D�4[H��{��>Y(8~���S�%0<7=�V
f�.k�$��0�H����ݹ1Zd'~n�F簧%�Jw�?�h�h�Ҕ;ߔB|��fc��s���G��u���	e#�gk�>���S��㾑�UFu"�&\�E��k���'�W�fk���sq��	��;s � _���Zm>#����������տ���.Q��fޑ�ee�|x�"ҍY���WO�b��fS���M��`SY�m����ʃ�pC�bi��8����&���!�)}�b�4ەt�Q��Wߚֽϯ�X���6�G�w��3�{ѓ^�|��jM�-�Ц�ږ�K�c�OK�?/Ee�z$�^+�(�͡a�&���t\j��$���+ۑ]d��2?��ĞƉ_��
�C�ɣ������}"WN|���⎃҅�Y,�H���W���.�����.�{��w��e7f:,�.��c���,1��Ԗ�ia*��h"�(�������co[�`��Ԥ�����0�qqLŴܠ�$�%r����İߦm}� ��ii��oo�E�q�𙢜t=���>�^b��{�{��[�Ns��c-�@������6���J���8�3Qk��Zbu��\ �=j�4ɭ�M�lg�Q��%7³��
�clR��D�-|������R�!�萧�758=�&k��h:0��CJ��b�G$Y'�;���@m�#�r�S�M NB�p�c_�,��e6��*���8�֪cEx��zDU����Cو�٭|ս�T�	��bɝ*�hI�i������#����9q����bN�f�ܬҧ�aA�&�����}TK������q�t������&�����N* ](�gB�?�zp!���������9�3A��y�ל�f�Ĉ��8�3�U�4�m���\Lc\cVZ��T0��2�^0��~�Z\N�b�,�v�hn[JА9��3Km�bs�3�v��n�7"~8�#�^��Sd��d|��ށ��wJ`�@Bg��Xa0/�\�+*TR���j���z����_h�m�4rڡ�
{��[~��tD���#��{�gR ��P	g�?���[�!<�Ҿ����x���^��$�11O1 J_��#ȤX�yk�Y��+�#�9�H���їK�!
�n�q�����-�pc�j~��<L�k�d��,4�h�]h�J�Ҿ�7�\9WI����҃9vR��^$���/�*"]�z���j�5zp6�E9 h�`!�D�C�~���W^5�ةJ�����9]��� b���č�=��"�^�Kf���"�Ů�W)��q����#-ʌ�O��[���XjA�Mns4_ �K����(�
����e�o��?�£`���n�z��%�x�3Ui[?5T'����eJ>"n@����B�?��A�4�8#��"��G�Y��k��JV��v3b$�#q͊��W��G.|yd�~���c>E:�s�؍��������m���7�5m@s��cmy�/�z¹z��� D�H�A�ژxDbQ0Xf�K,^c�Ws�q2`h�~�պ�V���"W)��i���`x	��UӨ��W[��1D�>�I;JQD8}���u����alT��)�X�w��u z֌`���F?B�%�<[/��e_ݥ&��K�HFsf�8�3}䄪��c܊�*�v�Ɛ��HF�d�yY��C���q[ɹD=�[ӹ6ԙa�f�8� �����#�|A�$�.�9ߝy���Mlx�x�d�ϑ:=�5(�7ׯ�tuv��-�QNǂ6�ŨY)X��H�e�N��7��'{����7O�O���sx�!TK��9�8�d�aYR���G3f�u����t�mӍ��L ��t)nc�ϒyc\�o�4YH�s^�lj�_�z6r翶'��,{-p��:P�T?
W�D�4I"��^�T��;��X��*2n�X�d�����!��Y�ZےL��Si����@�������o�CV�̪<֫[I\w��Pr͵!�̏�ݺ�g�t����{�0c��|ۤ��p�o�����TZ�E@�)�m���D�2HZr����z�VA�Ĭ���V��cl��4�����5]Ō?�J�;l�~G�����Q�h�+�#�ŀV9>�Sā"�(I��k�3y}SE[	ù�{V.\�Y�#�9pհ3jZ��������T'y]�������$����az��A;ک��fTjrX�0 J��2S���ʆ�7#3���I{�ֽ�5�L'	�mu��fA�翫��=�"_��PI��p~~����0 ?]J��3���o\S�����i��c����/Q1�Pr�0����Ҭ��qy:Dg#�|��֏@���Eg>�X8�GR�)�9�.�qA�,Fu���Cf+ն����4�r����]5	�ƓO��Bk#N@�Z����e������� A.��yhe��w֭c�>DF䗐;�%�H�^��W��/�&t�ʛ�"!3�����6r���ٲ��byS7�D��t�����'�����;�VP0¶6r��� Ҹ�����rL"*lf��?��#��uu2�J�e���o���o�@:\�:�B��l��$����#h49�b��(Ғ���J��
CX{D븩�0�Q�`(�9&Z��i&�-:����������H��f_b�-0���\�5:��S=�uQU���3V�S
��S41�/\�	�δ�����3��4`�i����~�I?qs�d
��ݕ��}l�L�$�.���^Tױ����<~|ח����>��Y�lrCa���	$�y^�s�@�	���=�\b* V)v�hc��+H-�	��	�0��4����/D=�� 5_�g;��։n��{��.��^Ȕ9�M����~$�]Uߞ"�$D4D|�:��h�QG*b�J�F��"ġsLw:��9�� k�C��C�;�HD��q�� N�P������/z,B�b��8���|6��:��G�	T�aVy�T&z����V]VҪ�r缐�;���hzl���8�����p�	A�a/��]v������T�6a�W�^��8	��t˯wg�h�[���1����u��_b������s�|!�b�!ov�V&'%���Y���&�j�s�U���i�]Hk���T����Fy,E�`�\��(�ϻ�\�S�<�*�e�-ʧ��74�=v�-��xy��4�ǽ�ƣ��D��W�b���j��[����h�SDu�s���FhB�7��N����E)�a�8(i�MOy�ei�Ѷ̤.$�!���\��
��d;�w7B�߽��F�����/��j�܇�����^�L������;�g5�i�Q"l'�zM��]	܄e ��x�$E���鍧<5�� �}M�&������#N����4��]��ܲ�`U������`���f���@[6��m��g�4!պ�]:?l+�!l��_�<�T��~UhI
PTZ��˿b�%FU���چ�ɾ�����Q�Nб���H���M�[�A�0�*�K!��ꗭo6���Z�ll��9u>�L��	�n:x������n'՗9�H�_kR����n�`M��E�`M��/U��^x�!葚�]B�6���������|�#��P��^�",��FH����k�XM��\a�b�Io.nX�B4/����B<.>�5��xR(�_9 ڭ�^��̭.�[q��,����>���KB���p��_/	���`o��@\�&_೬gʘ�����ow0����/�/��J��a(�*r���J-���i�y쇰��
��O�����8-Hc���s�Ik�j�f[Qʤ�`P	H���x���kBs� ���M�����MtGw>@Ow3�CT³�j�e�[e"���#�0=�2��Әl�`E�X�NI3'9�!��f�:p$��iE�C���U_��|:e��Ql��m��N���q���T���؃�oQ�)rDH��;z ����j�p@�g{�Mwۛ���Є�t	
����	v���O~Y��;��(8ψ����~�칵�~L�Eq����b>>^uE��fj��c��̵�E�31y�`�7��t�RA��sc������b�&��������
��
�F��Kkt�/儘�O���oA��;�p���݀�N��P�C(��7�5#2�%����7�&��R� 0�b��h:c�|p����g>�]��;=�����ۢ��P%�q<t�0 �[��Y,yµI!m���Y�ܤ|�IN���<*1��f,p�"���v*!|�����s�xG;{b�n���i� o�S�Ɉs���x�fO"f/ΔN}����}O1�?���Q3�$��Ӫk~2����^��Cr�ұe�jr���FZ��Ś��� O��5oO�n1����;Q&W�N�f��L m���d�7���]M���s�DZc�j��Mh [L������hWn���"{x{V�|�`���^"��+�ըs\�nח��y��bV�Dkyӫ�F����K���Fz�F�l��=��@�K��K�sڌ)��&�S<�g ����E��l155Cy���8�c��*Pk�|��E�խ�/N�'�Ki���.%ď��<K���6�� zHw�[��֙��D��ښgB*����}\`^�L�	n�F���q�=)��#gv��<1\{�ܜ�Z������{�I�f,�F���-��1��!q�U��S�����$�$�r��L�N�4���C�q����^Ɣ$ւ�Qti8�0O�+�/6���~�OD a��+�m��t�䷺�o�q�p��;��.�2���}��������&�(�[�v�qz&�t��
4C�t��񅀫�&CQ�^G-���>+����'�H���؅�\Z�SN��ymu�<RM��^�bѱ�K7�M�"D<6e��ƒa�%��m� ���ղ}$J�Z�%z�6��,Q,��vS�Z��Q�׷�&A�2?��Z\݌���KC����T�U���Gn�'_��䃐6vu��kOQW>+�TXV�s}�����TFnݴ/������V͓�>9I��m-U|E�h��3�
&���6�^�Un�9�}+�Ua�.g��h�e�(��o-�ֵ�k��-a<��������ݠ[KJ�I<�<Y��!�1��~�}	 �x���&)_��h� <��G�a�o�u�f�h��CQ���&0A�ۓl����m�����Iܚ�+��O ��=j۾T�	 �a�[)R�6_�K���_��/����5z������zq�yD�AY���l�\����T
��A��C�-I��t#@�������F�C�8	��w�a��<uo|���Ԓ�es�=i|;gT �l�3���	B*P�=���7�S��1~ ���ൟ��*�2�uo� �r~�-+�׫������R﬷�V�����^��3x��m�O����@�o#?��i�Ǿ�OϬHJ��9���u^�W����js��e�W�V�������xd�'�ܦ~Tӟ����`Ʒuo���$ Ҽ �/'�W�����F���娇�-G\1C�ՁK�bk���p�.t����窜#�.���^�Ÿ%_�G#[�#x�c=�Z�)��KI����^�,������Kr-!
������]�C���  �u�/Ŧ�?��F@ٞ����6%ᑴ$��A�I�b����P)q)%s�� s�4��2#�+ꬕkF��`���a��Tԉ�NH�3�P�x�(t��i���T���T�U�K��2����,SU����� J���u˭��q�mHl5g�������o�t�����.��ԇ�5�^x�Ť<{�n��)wZ5��#d.1Îp��f��Y��Y��zV2@�;W�]Q�OT0��W:�)�"� �A�^H���"����a�R�ͼ3~+����i���6��������6�A�;>��c�n��觼m��;�:����}��7a��6/�s���{�ډ��q'}\H~�{M~�TK��ŉ�r
��	���ۃ�H���g\J�Su�[�ȼݸmQ��\<)k��_K�\��'���U��?(��&V�W�e���V���ruB��_�jt��r�؝�������U0�f.�RSp�T�Dۋ��K�0�w��{�tD� -��;ϋ������
¤;� B_�ի���Nr;¿t�S��B�2:��Q&<�X�(����d���m�Ca哔�;둺F8ٖ8O�j�����2R��-�n�6ę���#�׭���O���&ԡ>hc����`�����Z����(�1��1�^yu�[�����D9C-v�-���
�ɘj�E�9�<W�7Z�T��j�ј����FS��I"��t�x���༠�b=�CM��G1�v�a4�(uj�N��KZ��ŵ�T�ӛ�2M@c�2+NuA�@�tn���!9
B��B |�[{A�լ-cJ(�$&�+Ϡ�
ް�	�=u�n�����7��	��J���U��6����ġ,(ԧ�p�Fhj��;U�`Y?[����d4�esL�ԯ+�2����V�D����}�ȡf���l�^�}���Y?xo�>�������=a�HK�<;�xݸ����gEtR�d d���ܳ.��d�,�{Ǔ��MP�����W����&\���p��ŲXdѤ|>���Ii�2d���S
���G;�f�����8bZ
p?�*+�rL�	���L1�EO��RbOqa� 7�:<�+^f��tw,�����79v��$�ȍ����εv�9)���@5�ۧC��$����7H�u�8��ŨA{�C a(r���0G݂h(+���dz-K��r��G�fq������!��
9~�������?L��:�����i�@&)�G�BNHb�\�pMԕ���x�id�Z�M0�E��Q�6���p�&���L��P½�q �FX��N:T1����C�a��n"}H*%6�`����m�~	 �#��M bn6<;��n�F��~�y���V�k|JF0�+;��c��F�V:� )Z2�bv=_V6�	 c���(�c��h�H���}��b��z��|�P%��o��&�RA�2��$��+#�d���Wxt�!����$�>P�#���m�U:��f�C��(;4��)�<�$��E�N�P���l��\Jb}���6M�D���� �֒�����F���J�p�^�Ɩa�i�\�u�-��M�a���vFv�Wsb�a⵫)����}G/5]��'�ֻ��w��Gɵ�u�w� ����.Ÿ��A��m+`�8�] V��Fi?�/]'�1�2����>S�cd����}dV[���r�)f��fD^6�I�����՟�I�&<q���l��������ȶo݌���b~��$���C\��E����k6vS��:�Ja�G*�FV1��G��Tj��6���иu�ܭ��J��/P\�3������c����(�P���� :���6E1Py�M�?�&xT��'A��4���% L4�{\D�ae:�.�V4���\Qa���]$s:j6�cXE�;t��\S�_W
�C��(��
����y��z����j�$�%Ju�	��/��ou9��S;-��u�ź�������S�g���7@�?z��xL	��ұ}s����$xL��E��8���xyp�����q]���e矎�n���L��+��@1<-�qǧ�~˅�C�g9֋&����YLd��	�ҧ*�@כ1�+rR�o�D�<�� ��1�7t;[u��*��Z�'��n!w1M:�w�v���D�Q؜M4��ӻ4��F-�u�ճ>�P���}d���ZzMY(D�|S�HX���1�o�۾�D����V�9�-�j������J5wh��@�
}����ȼ��ZwL&��n�|\�	����.��;�U�`�w:!u�ھ�2�÷�&G�&ET�϶OD��7�]�����(	�<�w�A�&'����m��|�T_ ��"�fmr4������LYbg]�9�����J-B��X"���_d��$,41oҡ`�-��m5����o(����+�6`�R���*V��k�P����)Ś7$Hk� ^D���
R������n��#��;��D�����?��0/�~�+�yC(��*|a��w�1��3H���F��F�S�3#,*$ؐ��K�is`�*��@\��b�3q�?,�%R����z���8~!z�7����u�>��o��9��T���g�ge�o��� �.H=bν%b*���JD)~����M��6���H�A��_v��6���ns�z�-0|��L�.��S��t�%����R���֍��t�W�7�dIt�jT���B�V�0���n�
�I�'��Y�nB��O��꣕��"�b����R��)�ȍJ�����Zc�:�I�\�2��e��qQ��M��2�Z"�5��G#�7�]٘[�ǢI��ˁ�	�e���e��}3C���{�I��o��d�>i2C�X��hW#�⥥E�
�[�{����cC�S�,��s��9�Y��F"�LE���M��gt���;z�����S� ��K�/��_�T]HV%�N��|�I=���g��4�����Z�W$B�f^k��#��kX�n��I\�K�q|���GSC7�!I1��\i9��iO_	v���[�{����z��(�H�k��GqC ���IHv�T9����{5��A�);8��Oy0���aY?ء�A�� 3B�m3�n��솤�7�\��!q���[���SG��A���@.-/�w�1����f��<��m�_�}�j���'FfT���*��KE$j�mu�m���m/�Ø������h��5�!�q��ğ����Y��"��Y9!����G`����w�"-Ch��ă���3�A���f$ZS����Z`�,=.ڀR�M���btLh��N��0�$�A��Th:�Tjz=����P�GH��Ӄ9⾑���$�眦/T�ho���%��KX* q6�-�6�����wU#����Ӡ�!��&+t��׬��uL�\x HLW� 7��.'m��;Tݔ�c�=� ���dn$:� ~"q����{��f|�g֫R ����d�O��ԣ#��l��h�|,�M������rb)����]�bq��ȇLW��WV�>E.��FɃg�v<�:a�p,jP�)|���6-T�|$G��=�]�o�,,����.�@,��ʨ�~�k��w�TW~��ۻc�#��uFbyŶ�y�ޱOW��������:�nݽ��p,�R���+߅�_ �����{q���(=Bf���]��_A4���Įt�Y2��݊Sef��_H[2 .�^?�g$y����F�䇕
�i�@ˋB�DK�`���U��&M������s´�R��p?����X:�v1+�qV��2�P��6:�,%!�1Šm�e��2#�^� � ��mG4s�iX��Zm��N�<Y��`�1�Ds}
S�ꅱv�9lE���	;�Rr<3u��%2H֍6�ǚ�0q��Q�:Ҙ�6dܘ �m���nE���N˽b�S|�:s�꣕r��h�C]8B�r��Q�mZ����|������"K��l��_H��4�5�J�W�0b���wb�s)LY4:�*�����4<Lr���'}����f�ؕ��[]o������.V��o�ή!R{�Q��:��
��Ke�Gh�K�;o�����*K�t�{p��Go�#�a5g���\�������|&8�ö;/��J��xt-�zTF5�
����6?i`L�������$ �WxX�@�/��(Z:���ImF�2����_�|q�`3�"���4�46�����/����q3ɾ55s��b�6����.���;(�����1-�(�F�#n�7����Hw�+B*:76��@����_mj�}IA��r�`$ė�!���O�R킟�5\(#r��a ��1(�]8�/��*���J�O�����m^�-n�����f�z�x�x��vZ��"�\@25�3��K}��E�p�8�\c�%Ƽ�c�Pʇ(E�K�b���"�P��{c]0�ok	ohp���Q���b������il��b�ԝ�;W�y?F�g�Ao�@��r�J�~s0:p-��#�9#z��&ٴ3�9ۍ�n�{��צ�j,<�I,�G�i��h�#X�2�5�jOBr�k����=�#�X�Z��a}��x
�"����O%d���X��~�����:}'��Rˀ�* _7SdEe��6���_Zeu�׻�������T3�r��ͻ{��D�C�dsY�^|�$4���`3��Ca���0�������F�'�TN���H��߾Ŧy	vE;�q|�/Ό�dO3��E�.Vu$GJ؃�J�]4
T/�l4���Z��E	i a��L��G��[D���,~i�)����	K(cB?,1�&V0v`�+��$~���Q��sS$��`�Y�W��,3v���g�C���t�.�6�Sɥ�g��1�ڲFjj��ď���8����/h���"~�@@� �'�����v�W�~���evqhP�|TX����p}��,��L��e�A,�'�EbM_Н-i���C)����(]E�ÿ��%Di�TԤ�S���7u��OŦv�(�҄�tE�S�j���c(�����\�;�?qӷS�9!\Ryn�+x��	�n���
!�z�B�f�R>/��*}�Vˠn�# q�I#���n%{��������Ǵ�<�}���ďh���$g)VAr��l�2��E���Do����V�a�E�3��_�]v!6Pؗi@�4m��q_�~��B���P�jR 0g[¢��Ȉ=*�O����-U���He0����|A
-W�ΉU�bzy��-H�l-F�a>n����,�ɼ��ތ�b�������z0~�E��q��&�(7İ�Q��w׉�a�P{p�}����j6�����PQ���;,��*���'ɍ�@��ت$w�+�QZ,ӽ;D�	~�H���÷���P�[F��5ڡ��p�������n��B�Q�J�	OxTYw�d1�-�٧����O�~}�ͩ4eNnv�B��ӱ�Dն����:��E��N᜴���[���Rk��	*���Cїc�_,`C�J�ZWn�k|���z�ɉ�خ/g[�Y��� ���!�+�rK���}�j@��H�.��T\��ލ�B���dfL��ivƩ�=�w��E3i������&`����6�,��rfm$]I�ɔ���Iߋ)[�E����ހ�r�Pl(8�M`�P�B��,�w��QXU�+ϙ@t�����^y����/��{4�����2
��06L�k���o=h��ԏ�yz�"�c�=-�XM݆^�<��<�ނ�L���(۷G(
�zwq#I��$�")���[��:+�t��_W��rj �t�`��^O�E��q�xyנ�=�i��SW:����[�z�$'�`=_Z"�w��E�i҃鏬��)�~��rZ�����_0�OO8%#���@@1f1�*]w%�߂+��.	:P���&}E��~*�����iTx)ys��ܐ�T2)��b=�o"�jϬ�'�C��-^���B�esf�f'f�$L紁��M;�E�u(&A���3F��ح�r���*X�X�j3�\ϝ
�{Y�N�$�P�u�Hv�z� A��4�\���[_�̷1�ʏa�Xгm1��$�e��{ɇ$��˾���Bj�����b�Сv��cL4X��T#O�0a�b̒�&|o4�I�����a�>�������Ɗ�ޣ���r��uVS)�)�N���q�$�!�5y�$�Pb���eD�8�uT�
��~2�/)��>Z����gθ"����C�3�;�[��������-��uC:y����r�����e7|��)#�Päy��t� �nE��;Bg�)�7��%�����Y��P��b��h�rb�F�sx�'��g������Z�:�܏��8Dդ."��9�Obεx�,�*��e5R��&�U�K*�wv��X��Y�a�4����q�kB�4���9��
���=4STy�f�����df|`�`��_����Z�����%l�Y݆
ilN@���עw��C�O�~��Vm���AÍʟ/-����=��#�w#7����E�;x��\������k�8��	�*��Q]�uJ���n�H�>� p|$(�M��T��m1�Gw�a�"����P<�ڃ�&J�����Vz�Լ���h�>R��Ps�qB�ҺX���L��!2SE�4{�A��E�m5�%�<���2Z�Υp�k�hd����!;�Z\-���
��=G�geqfߤ��5	�˖xY��"�]��87�'���������w�z�IO������%�%Y� ��%�8���!ef���`����f)t2�#ߡ����rjXnH�C��؇�eǍgqz����.z�0�ӟv�J	�+���U��;�{����g:S��ݝY=��F'6<Fq�W�.A����ycm`�z)�,���ƪZ�o��V�j�~CYgG�Mc������D8��m��WU7U����ewS�Z��?[��m��� �cˇ	���J���v=Ҕ4��a(�A���%.�X�H��-�kt������=�%LʓC耎�ӵڥs��Z��Z�KoX��h�hY6	�a�"6�/ɾt��٢�6�~��oul�P����$IfR���ߊ�7��	/3���#�m4 �Mg'5=��n�Kw]6U�FA��:fTt�+�,��khO)Ŗ�^i�+�����hGp�D�]ay>	f��ݭK���i�qs�q�߫�1l�|��3��L&�`N_�g~-Y���AN�	j^H���n!S�k'T<H�@fP��]R~#^�#^z"�"��0�٧��G6V~D�C��c�Es4Ϛ��Z��R���
~���0a�uqسT����y�'� Bˊ��߅g1��sh�B�Ȗ�]F�o:P���b<���C����1.P���ޔ��Q%b��bt|��.7�\�i���$��نx��"���d��%�3�zc<�Hx�<l�k�u�Ca��Gt�jd��c��TY�om�ҏ���τmhʡ��d9U�u	�s�X�e����聈��7���^�ѫ~�g��<r�3&��;4��M������C�����3c{1E�B;�Hv��E��d,�ah9�.�+��Pm��~�� �箵���rTaʣ�Og�
�u{߉��!�G����=5����Qkժ�g$�[d����c�Y �����?Kf6s���ÿ$�0�|�i�Nͺ
��)����q���X���V4��c��2�}���Rwf���I���е�����w<5ݜ�d�#\a�w���	�	��
TOO��/���2�(��Vb�����QΊ�	UC�d��qkO,6�G��3�kҘj���cH!s�l�H\�y����@�t�zq���BF*ɝD���Mu��7|��*�1�U:��ߑ����~���)W-6��G˝ 7 j��١����"h���sH��/�+>'#��	�^�1^NO<g d�A^�1,����K5J ��;ݙN|Hh]�]y�� Jt�Sm��n�:f��̣u�m<�V}L�E�E�#��@LY��� ��tQ1V�5S�;���d�+��4��I:'�[�F��:Nj�[R��-�K�򧡏%Ǔp�i��֧��7f�Ԯi�\�S쫀�~�����zH�P�)/�$s�Z�1Q�0f:Y
����|Uܓ�d�K�� ���Gw���խa�w �a'���X`Z�S0�Y8���ϔ����V�ywb�s���Zqs�㮛�u�a�GWmYh� _M0v����x�[��SWkX>uz
KG�hsY�G�N�����	���t����4�&ơ�c$�1�{�3:���̂��� ��1m-Qf>͘K���w���#V��pP.��e�s���yr�+�T~�Kҽ@�O����.H٢)1��0H`C�ɚ����,�
{��#���a�ao�M��hx�y��`���B�=_:ۏ��O>+��0(����cX�-�Py8�s���V��S�̝Dy�Z�#��B(;D���8/S�*�=�Y���!8o�k���*)���b�z������ͮ.����Kݗ�˻���
,V���V�y����7Wԯ�`����	�x����Bʳ���AtZ��`�J�-tߘ��Lr�o�j�-s�����9�(Z�-ۉ�=���EL1�e:�������1�NU���*|�89��#����V�BN��J��O��F��m�Q�D{��h���a���\�]ʣ(ފD��D��TdLGĨ'�G�oVV�Ÿ�����܂؅�RB�z�m�J�_�H�M?��}�)��M肗�^nY��2��	�����&!����zpK����<e�zz3�pBt���,\���ܝ�����xFC��@y��
T�[���#���(i�X��g�@A���x"i�*�@�yO$��0��&p�Ô�`��2v�6[ߺ�'�7���e�X�!P�T��D;���/�[��o����Dd��x��P;wƒ�V�,0�YV�Nq����H�;�E��m�?�O8��=���.�x��(�N��{��Qw/?��,��UOS>�f�Rg���>��(�� DłIm{q���@���1�2����%�������Q�q�ח�����Z�E�9�ǈ��	5
:���7���lU���i}X;I6Bj�O?Q�	<��~%���q�X����{��B�?^��3Ga���ȾШGM���=$-�G�9�Q���8�_"&�ҡ�=e����>J"��cI��s���,IQ���1���]C�^�?4�X�]Ʋwl�j��8��ʇN�-m`�7���2��/G�=)�ɏ8�gx�w���t�a�����|�(��tg�c�%f�
X_���|�0Yv���s�6�Ä��Q���ݿL�H�X��:>v@�r��;�f���}���!~�ھҷZ@Vp��j�6o���c?橑V�Հʝ�2 ��(y��O��8�j���!�|͵W�2�5=ԥ�d1#Dy�3L.�ﬕ���3���e��t�g�#����˸8}�Ǧ����+b�����j�\Q�'	��5���'HHO���������6匘��������ic�HD�� LNei����}bV�(���Ԛ���-f
`��e�K�kO�����쟅���$q�I����5[�jJ�GMF8�̳���W�6-��8N��~�8�-Mi�Y�
^Z�-s��x5ù�u���vA�����Z��aM���F��v+�����o�̶K�ڀAq��%C��	#���
%�����TK��U�*aE:�܅^Ec��ڃ��۬hԏ����xL�"w�w��Eh�b^����6���6�t�p���ȥgF4�B�g�	������5��,�̴���������ѳ��]���%�U��OLe��lQ�|�~�F�{�v\��9��ځ
���x���w�i�2p����4F;�f<��@ׁ�ν��w�#��uh�P�v�{k�RZ��������/�W�a?��m�Dg�|��V��	F�T(
�I;o�S����T�0�Nr��	36'Ӂ@�(ppo�����
r�h�`��+�m����"${y��	�]������⬚?�����ծ9\��'�X��!������1�v]s��
�����|�ePa�����u`��yN�\��Nl_r^������N\ �R�쳟\b�@�"��Ό�
�hY��3\rF^������//w
���$,O� zA���s|wJ)HZ���x~�}�4�ͅ�=�7���.SD9D��?���@�MǛ%S��Aح�~8������p%�"췖b���1�1���Ϙy��ڗ[MGV�h�(IV6'!x* },`�߲�#��� �1��9]9�3bI�ҩ��2�(?/�iF56��������1fO�Z�2C�@����=�2�uBH[��C��������JY"	j65r����eN�*�%�B�W�p"R����%��<�{�1���X�2�_;��k���υ�#���7�|�^_�X{� ��i��I�*����9�D�3�Ĭ�A��nd�܎��D1"O��<��.�/z��&90 P���m��E1J#h�1��챕ΡG�:f.?�l�� I>�?�9���[��MSgF��58cX��N�t1".����'�Ed���w"G�������2nҼ9˗�V��`��#g��I_L;LM|,d�X\"@7g�mϡ��4�߸b���B�^/���|���RB^�,M"��E���/����>��t-9��q��Ed<�G�<��P⢩Y���$�i.�k�+�_Fy������Si��TL۶ɞ0>)�i(?N�<�G���O��Lu O9��H��:��r����g��p���q��H}�]��⮛J��k"X�ؤ�8ճ�fz�v���5&=ȫS�>X���5:D� �7j�0��ׄ?57�h��#e�(���wV4`lU���=s�m�Z"K��YҬА�B>�����>0U���4!Æ�L��q��:WNV.� �S�8'��|Nd����c��Ǫ���*`��#c=�2�k�D�m1��y����0)�:s[D�A�\�e��S5�Ϣ_Y;�q&Ф��U]OŪ������`-S� �m�⇵y���M�o;?!c���=#�k2��k��A��B��%)D���s��2�3��AV�mO7{��!��<&�����<��^�O�[4/#ִeG�I��l���f��EqF��5�gY��Nj��VO1ˑ�◣���7��	<�.t�,怤x�&EF.��ٽ�0�#���
����u�-����<lD�&��E��1I=��@��a[����i����G��`����D��9e���OK���70̙���9	�fGc�w0���>ѰV8J0A-�8��$��(�$zR�`H͵���8�-��X��i�v;5`Z��Q�O@tߐ���-���>�9Z��ub�TA;������w�G�a֨[�����t�)��ý̳���L����Ḵ� �b�nu۫�##�u�O�/ˠ��͎3ۮ`T`M"W�<FB�6ö\}�!	�Qc��� �*�?��=8�`k�l3L+����N�a�~�+0���<�2?�VJ(�����yĕq��.-��}I�L���,vb�p��k)ʐ�^�M2����'��ލ�O�2f���m�m���ZŬ�����,�6��1�Y3k����<~F���+c���`x�����a^�#��/�h��_��'fL�iì���gے.�nH1b�n�ߐ1�q���'�AƵ�]�>o���?̋����5M�O_���[��q45SHXm��H��������i���T�#kp؍ϯ ��`�m��i�����zJ�u����Ӛέ�.Y��� $��?Ѝ�R�|�( R��Ƹ3�z�c�0:z�$�DZ��n�[{W\p9��N�p��@9��5��&f���^��)+|DH��Gb��N�]��F�o�B�0�E�!�,�ԁx��3�
?R��Y����ry��O�9#�:Ɂ��rl:K%�8��jd5VŨ̗��"[|�.xm|ş	��	v9���y}B0:i��X��c���8"x*7E�Z�^�VT��M���'e�.�3g�%��B�ٝ:��<^���_�;垪8:F6�A!����m�����9�HS,�r�נ�gwX�n榳�bq�kc����L;Z\ �	�I^A�s�i�p�-�7P��ر����Y�)���e`�Ǭ$A�ȬF^�����#Y>��)�V�Ҕ�F�fL���
�����i�ݿI?Ҋ�7wE������ٛ��}�i�h�SĿc@�J��a	��76�Ǘ���,!9y��8��̿`��ȊZ5$��캋z��n\���ɮGB=��m�Q�m?�����Gd��Ϡ���ᷠ�_������'eK}7D{<��H��R�7CVR[Y�c8�����������v��x�������o��	y��iQ�+�oSܑj�����[}�-wu�x �����;j ]p�`*����u��B�� ~��.��.ވw�.\���k]4�4d9x_��{��<���T�Q\��&^'�ףrc��3z8��y���%�}{��f�t����������9�_G����A#��{�t�iƅ@In�W����-�@�ȯ���GF.���rۤ>ĉ8��K�)'l��z@Z��ўӞ+Y*�:��L��݂�Hk����&R�%���Pr������ht�!����FF9�%!�P�r�;ŉ�C�p0SlS��������x���g�/X�����x@���|�@�RK�j�"�Tx2)d,��N�u�$/�*F,�m]H �����o�.b��LV��r4T	a�Q�d�z�P<�p�[4ixq
�K}tw_��0�B���?�NLǉלU�o�u�"6ӏ�*.#��z���g�t�~�j;/�M^K��4w\���dj��iL�9]615�f�:�)�\z�~*n,�&
�~���/�\�J����0y-j�=�ݤ�Ӱ�{��,-~�_:�2��d��
��oQ�p�yb�� ��:�s���Z]8��̲�)� ����n$�2�<C�S�Aс��7}�G�����F��
i6�G)��x�
���^]�o��q�������`����
���%o�����r����0�][��� �[���� �q�]���o5��YQ��]���l�>���NfBn��ܾ��OT�u�o��Q�&6_�H9O�Ԏ��XR�}6B���u˱s�$��������S�[z�L��l��]�}כ�Kn
���8�N^��M]�Ly�e�}�U6R��UzRh��ߠ�Wr��� �����1S*�D��B7������b%�#���@�+�bS�=R�B��*35=�9_��z�� �����=un�^���V��BWƬ�>S�T|��G�~l��T��}��H�]��^M�
��JE�'�=ƙ!��f��'�H�U�[�E��hL��EP8ڔ5��<���0��e�j�:m��a�{(w����ރ.��	�-m����W���2�� �!]�w�z��2�i*��X4:݆՘�S�E�#��� ���ԝ�H%�U��+�T�0�_(����}'^M2�h>��e�[Z%����� �O���|�P�-���ɖ@�;N��}1���4"F�ǟ��_ԏ)�d΃�EJT�d�p�n.�b�ƤɄïX����_�P|]02ET�N|��G_�FPnb��_�IE1E`��{_�׵�.^�/f ��n�8|�2S�X�X��d-O�p�����n|�Cc�6��aIߊ����k�\��x�����9�NW仑��|��降�8��YÑ	'�g|I��n4��"_�0>�!OIUi4`gY�a�5�	���vCڈi�x>S�	w4���ԽrK9C�X1InY�h�t:�I�)
g�w�qP��Y���Z���R�"��`F�4�Ҭ�L���V�݄ I_F��qlgӰ�H|��"�A�e��ܫ�����I�� b��O�Ti�H>N��`FS��Y1z�n`y�m� b�&�{���Gc� �,����6g'79A��KD�����FiM_�er/(a�iqS6�&!�h6��\/�fЮ���
a�nT[F�׍߽�u��\�A��ݠk��#�*��9�b��΄��g�U;80�ø+mX��M�z�BI���TG���������@�����`:܏��2EF���t�;*�_�2M~ZgO�)�M�a�\lС�4�2³nH���ca�jE���?��p����Q4Zw�W��u��}M/sl\�-��z��'��/���@<���LMK}����B?�.#���h�,m7qH��E��H����7X͇$�=	����CU�2���M���1�X�^^�ʅCHJ³R`S�~o�Do	߻%L=+�:ȿ �x���R8AX�>�_f23iaO��������g���`k�if�/i'jh�a%���\�����-=�&���~T�Xz����!�����7�aKm�͉v����}�BDzP.�
��6���B�&8�Q��	��f���DW��vc�����~Vb{H�c�_�T�<��ʃ
L�آXZ��o�Z/��.��U��@NJ�	��QB��s��+{T�j���R��'T��e�%{F	
~%��(�K*�j�Tc�v�*G0��`��������&M:���,˴�U37Љ]��bO�8|�W0f*�>��q�̘~�	q�҅�ӎݬ�E�M��\I�<�*�fᕗY�o�a�:њ<m�������\ �����,��u�rM�E6�7�w!4�@9�r>�@V��0�ɦ�/�XN#���n*	49�IZM�=��j¶S���1pI��9�p�6��J��Δ�d"�\��wzm�B�Ҍ�0�|_ҮP��Ӄn��$�M%�1�E�^��/�2�Ȧ��㴴�.�~]J`!�^!^��
����LOj�&/�{��Zt��������޳� �����*����}�_+���I����q�x�R	�痽�`a�jo��������%k���*��~}��W?��~��y��\aM��`�(	2:#�Ï�g���o{:2xg"cJ*0��J0�%rmM��;��/���Dpc�eİ"H���ʽͷ1/�>����JU^��M@m,9,剶X���3���cs�t�O����2�����W��M��2E*N���4�v�X��_�-�C�¬i��NG����h��EU,^���m\��&W��� �e����t\��1,P�d�Fs�� w$K�E��3X<B�(8��n<ؤ�P��ZB��u���։!�H���j���M�!b"٤d�j(��ir�d
�i}�O����-�Z1�B}�B!ϭYշ�k}�\�A���٠�T�<���~����$��(�j:�Mf�;�q�i��T����P��Ҕ6qy݁]F}0�O;���;�CLl6#�Rk��z�5l�6�/�5��F�io�m_�^ԑ��S�$!��Z�n�-�T��$���� �F�!JL��-P�sӠllAm�ꃸ��X<�e�	j2��{T��>R�<cAy�v���:&rN��A&�CL�/�9H�,.���g��S��H��c���Ȗ���T��ҵ�ZUۻ��R.�Y��YmA���X���mԃQ�bI�����r�G�n^�&XN�?�Ɨ�nS���@��n:7Z���RlՒ���sa�`<�!1~:O_��q���|�@v���`��������"�]�vwE����ܬ�Қ!e-���� 6���9��s9Â 6���C�����wk�v䝇W(Ę$#���bů}���Lq�r�W�kI��x�'���3#p�f�T�O����P$���	�u�+Qp�n�$�ZHJ;w��Z����3
u?T�����I�y�rw_����;/?!H��'v��<���:^$޵;tH��Ȳ�UO���� ��Z�rџ�T �Hp�<�������)p�y��Ԅ�V	C�u[��q�V�#�jJ?�#a�).��&@��3�5��� ��?܄�R�Z&l������?P�QVa�y6��t�@J��XsB���,�T�� W�@���k�^`���m]=1�"�?�Iˊ'\�ut�b��Tz�Ch�����U���:,���^*aY�e��PW|<:��6۫��a�{���N�mdd�1�D'�M�x��<=��@�Xa���>pJ�I�0/��jKxW勍j��J��IYBB_D���-�A�͑��Ks��<T�7�p�:dJ>8��L?������
��/ݵ4���H��H�Pɠ7�p;$�8�⊲������G�_���J��4��
'xB	^��9�N#��1y�O�*;�����k�V`5Y�f������	���=����l6S�7�6�lԘ�V�(�S^�mܻ���\6��~~N�lubI�d��H�Z�J��������r��%Hiy�]l��j�μ����'��&G��{�r���8jՍ��a��.Q,���w��.4fǭl�]j�C��n��&)ځ�.�\}�.�g*�.�9-2-���]ԓd�rT�8����?���l�~=&>
��� �����sP���^�P_X�Գx�������v�6B���X���e[�w'�GJ�V��A�&�&^�̜}��A+bI������5I{tyH5���3��i�Q;�h�`S[[cf�����Ƽ��5�lU`�x4��������-�kX����q�-��I��K~yR�Х]�G�#7���6!�;b�b�Z_��=6m��H�y�+�+�e��~�U.���΀�� ��]��N�:�-��.�� �=�*Z��1E<e�i��	��cDJ�l(�C(�Ò��R^��g6Y�Ajw�l w����o��P� �;��h�*ЈS=�\^'֥��g!���J?�dm�(C+�p�6��R2����r�{u��y��zx�D�GhʼB���������(��^�L`�E�Z�i�� �ԓf͊v.�m�ӘQK���~��ʉ
�$�K7V����{>h�cb!��+�!.�����������W��ab��C!��?���0U.��>{~���7�5}��	�P�u�I�J��/�?C
��ଅ��1�Q���*9z_�N�� ��2B�T��5���nH.�h�t���̅�&��׺�r���OY�k�Ѷ�V���,�`�7�*8�F;�_r�q�F�,��Էr���`�P���dP�����`|TH�OTŸx�#�������3��1$��yf7K��Ƙ	�@������8���p���sW�	�i��B���+l��N�ٸ��Z2���㱳!_5�VQM�z�TN���w|�i����H7}��4��q��B�(vp��Z�D1�;��9"7��=*�to%���I�(�/��DMp	̀AϺ�_���E��\��wg�HMl;�)"ǩ�����4�mE�gK�r">��Y��٭5k�h����?h����$�+�.7���mu�;�ƚ���Ҿn��2��+�#K�7��S��Z4o�mN��=4��7{���L�
�3ra)���"��8BK�?L6ѯMC�ـ2�_FP�0���O��qj��o�R�l�}|]�vd&,�0�nś,�:\�5��ؗw �/q��:v6���U��ˏ�%:�^ތbfg}��B��:~!(�P䂮�( �8�ǜ����T*{Z�h���g0e�����E ���	��4X{4���D}���B������$��"� [�Vb����]#v�ۢ�	���'�􎴩9Q�-�U��O��P?�.�n�Aز��r(��Ԙ��Jv�7U�C��Bg��6)�?�s9�ƹ�K}�!.���U���d�JށL-���=vʲ�$5(p6V�t�7��,�dW�Y$���oG������Ęr�`���SØ��9K�X�=�#�Ķ���Y��+B���S�p
�
�.����uW��B՟)�a[�����j�S�rfU&B[�-x��Ϭ�qQ%�W���x&�.)�m�0��?�eq����5	Q�`���}>"�ȍ�&^�*�GRX��	�$|�Ìga��7.#���U	�Oڴ�9K���`Hޡ���ڗ�u5璇�[��@lG���&|��݈�5Y��o$��*E�p̎���#h�?�i]/��G�9��0�	-Ja�F�=]nr� zT�@��S<���`10�/WI�hv�,5{�Q�Ӓ>X�i��2W����kYb�0[�����׆�.m��8O��?�	�q��R�4�&�~��}RFf`ϥ[|���kn�l8Ъ+3���'�H���ԥt��b��O��څ�+0;"�@�/L�Q�v�r��G��3g$��ؙCS��\�{��+�Ejڧ�;�=�(n�s�p���jEg�N�SS�|��|��a#���ĕ��x�:�UN�-$~��^z�6fm����A��8�#>�	� $?����"�!�̹��:-��$�l��-�{^s�H�&g���w�"�S�CkϬ����M����L�LD�Ȳ���$�Us>_�C(�аPvJ<��x�{C��F��*DR5��]!�D�w��e��xK.��:.�5!o&����'��]�ym��¶��`�� "�~6�@tZ ��j%W�;Ӻ��̣�ŧ~B�isU��L��D�`�C���	'��y���	LVaz �pK�$��B'�â? Y�wzNH�����x���taU`�khOhK�/D���7���&�ɞ���jě���(T��#�[tj�>���=Xc�.�;��Htk�.~�4��R� ��43�@3�*ND�_`.�Vc�����n�KyM����ҶDUf<����o��n�i�T��z�Z�ݳ7�z��ɯ���]ⵓx3��2�Dw?�I�5.?R^v4��2[����4�7I.+j�	x ��G��&�#!�8S�o���}v@x˳4�@��)B��C�*���l����vN�Wg�y�����wЌ���6D�]�_z�c�����l%��vN�Y��d1�gQo���tO8a��[VE����L�6��?��e)!��j.�\���\�����2'�y��Ys���e��qY�F���`���Fh7�M�F�Z���+����9y���H,QV�D�8�]��J�?j�l�=@��?�?��ю@���2��t@C�����z�̄=�g�L'1[]Aj��\�q�}�?l���=�\?m��@C�ВY�n���B�����܋��,V�t�i�5�hӷ�R${��$h�a��v�b1�l�XC�d�m���j_��"R���/jZ��G=x��ţ2{��z�)�/Q椭n6��.LY�j���X�0��6m�R��A�|Te����֛-gu��#ܐ�b��t���MҼ��:]7�y�?�hG"����b���Yjq>�dC���/L'��<��5��G��-YJWSӃ�c��>�X�.�ҧ��yr� ��^�i����|O��ygӛ�,�D� ۧ�s��1r�G�4rX%ˁaAְR���_pms��gZ�#�"�cd*'~�sg��%�8 U��ِ
Ȃ
%���c�k6��1��]��nFKI=��,����� ������%����;ܗ���L
Q�@��] �l)R�râq �c�G��0�<Nv@ocX����C�����]�it ���'�Gё�'X�߳�W�zt��]>2D�ZRP��� ��Em�u�[8*����ŭߦ��o�)�8غ��P�օ��y��� +�'��ޜ/bA��ǠUe�o�;� ����Q�&V���ŴT�����������@lK�DI�(Gb�������b�XHCF���'z8?�E��rU�t��-c�a⬑�1����fm�0!?� l�k��`�#:p�ܣ3��G���Q\ߪ|9�Jk���pId����G�k��dr�"�%�}�����ҽ����%Ca#�k2 =%'� �d�~�f3��f�܆�kI㟙~eڹ�.�dۇfJ�b��>��a�3�G���[N�͇f�׆����ϭ��s�-�`��;�%�Ƿ��,���n�?q���©�A}�+�{�z{>$��w���� ��)�
Y��4�� ���ע�0����&l%�����C�N�-Citn�/0�(vYxo&�{�m{n�n�'n��m@�O�W��T2�����g$�&Xz�S��;q���.�_R�C'�9�V�$�	w3)Y<�R��ھ}���|Ә��W��.5 �L�'����Q���!�'F���7t�H�!B����B��C���h�ұ��	�8�����̧o���޻���	h�(�����#�:�7�jD�<x���[KwM��Kh�-�B ���54� ���Q7��jGV�@E=��l	�<ҶG���W�S���~���%�5>/��Ĝ�4�i8��o)�e���(;��0�D��p���Z�[�4�k�)�NxJ�N<i���x'��=c��]�X�J��+�����	F�ނ�~�h�C��筫g:�В+P�.��r�$�q�S ����O�;�D�|5���YV7/��Y�"�.a��wԅ*\g|�H�y�VU��q��G�iR�'�g���V[�u�/�Q6r<`3	�4�;�I�l��ƒ�ޑ��V���Kx�rQ�il;�1��Lq��yvEJ�?m�
ko�#�3!���?v�Π�Mƾ��#JZ�@v�S�;�v�1iڍI%�sc���#�5(���y�x`�,� Fs��ѐ��ѻ�-7�"*�k�����D�l��>�r�E����0j��t�s�A�
����B�MK+D�v���3�:����kµ���P���=y�^Y.���A5w�5���汽��pj#��&vR�j��b�@� ј�������b�јchk� �4����������i��\�U�:�m�z^0�Λ����FH�/x����$+�8����9���6�o����vw�=0A>V=nrS"(!uȺ��}Gu�~�#j��{�S�r��o�[Qz��6� [zV�:�6��>^5�Jy�KtG[^6��_å�N����g�h�T���"�5���,�'��p�s�mR���U�e��8��=Z��y� #�e�?�ͅB_��?ӹ?�T�GԵ�#��7+p������h��$6��Rp>ލl{K_	��&�n@���W��'K���8>��a�Ჩ�~Fr@8`�q��ȍ�#�W͏ 6�(��x�����け-$g���S�2U��^$�i��ک%Q���'�"Tt�(����%�J:���,�A��c��?-F�r��lx���W���7#�D�sb��̮�+-_���$�>��[�F��aGrj�4/w&��$O��X ?2v�h��*q~Ƒχ����{�����Kg4�8{gb������ �P�0���J[9��¥"�]J��LƼ.^�+RC[��ܡ�ٙ��@��ڬ��VX��b�뤆Ɍ��`�K��,A$6��@i���'��4RM=�bŽ0�{/19��k�լd�Qۡ�&�S�(�J�i���p��������i{<{Ω!��&ޣ�	�Ft�@�Y'uA	V���D�o�{:�r���}HX����i����[�����X:3��`4J4Bv�*�0��MG���?%�WhP�Y"Jkcjŋr'�o�uwn����7�PRS�8gZƲ��W�'K&�O�4s��SZ�z�̵�v~��6���%Z�6"ć��,+�2:�I��S*���>��t�QB�45��ȕËϢ�3Du,ٻ�h(�c��P��1=����w��@9����2�n�uX:O�R�J))�e�9��l&���N�,�[�w���^r�Ax�k@�V��x�01$[
�����k��:02�J�i!��������a[E�T�xZ�+Y�d�:����e�^�����M�JZ�x��=x�?���6�C�f�m���g$ee�#=����-��'1AՇ��4]E��1#/�?2���JŤ}ߤ��åt�T�acp|9�O���rLm�����Жz�b(���q�T��"���w��wmL��n.�+�A�U:�_�?.�($o��H��öRg⇤��u�ƣ�	�~��:�g����L �V��:�$j�ꨯ"F	�
�Ľ��M}�U�Pwh��c.���N�������F�S)�Hx���S2�4o�z3�j��Ld���MV�,��7�NgP$ybbJ+`��'�@�`��b��ky@��}��E�����IZʋս��>��7Cb(���*W)Q�=:��8i��sGby�W�b� ܕ(��\�Y��e���L�.Qe��ү��y�S�nt��G�랼G*ϫ�[��Ckf�1M�2[�����"`W�ITU���e��wd���ի��I�w�]�c�#��|;�a5��mD"��v����J��u�7���B2�ځ��
��E�X�FJ�M���n5_`�5piXV2���g�6��(�L��I���^+�I�e�u���e�>|)�G$��|@�W��r1�[���q�o�i�lWF-K8�iF� ��Z^Qe��y�����YA8�C(5A%n��2�+��2���$�F�����#$ Fu&��?.V�n`z�悼X��)�!�_f'8�����}�;�����P쵣��ʞ�]5�i��ࣴj��-��b?,�e�X/��Wiߣ���I�Vz�w���&&�����x��ƺ�C߇��.�ס�����j�i�EaP� ��F��$�tD�vQ�vG�/X$�,���B{�j����zrܯi��3ݝ��x:ě��qu6���r	QZq [�L�0x������e�g(��=�o��
���ðS��N{�k�e��<�OT���!n��ͭ^+���%5	z)IBV���h׸+����
��gx���3Җnx�ݫSJ@u��}fťhjHoҀ��V�ls;K赞�PjHfi��Zԍ�bs�̉�cC7���"��i���k�|>��Ubrۘ8���T
��*wr���sw��7�G|���,���lŧ�gE��e�W��#���<13et�[Y�7aҼ��%th�~	�ז
9 ����ܹ����2b��4���f�}q��ߎ]��*W���ƚ�l������;�:�{��r��UB��.�q���g��ñ����
�o�rf��8�q:~i�0���^�E<b���I���*S%j��J�?,#IK�����G��.�r���M�l�g�]_k���_L�ß>P��Wm����H���򔗬O똼8�����E�`�ј��F���Ly�-���Ο��l��;�I�>.�g�qn����F;�Z�W��8�ֺgv*��TA�,z�#���	a�m�^tYIf��.-ݜ�����iX!��̪�����]�DP;E���H�y��9��C�$���/U��(��������rq|�@Ѧ�^�ia�&�1 ��yI���R�I�dh����o_�u"+�D�<��-�^#����Ow^�{jl
�k��ڽY����Y�w�R���:m���N��`S8�b"�#�ɿ���D�|L��H�M�J�r2`%��*���B�'�&�|#��t@d�&���[_�JEs��A�h.�H��ã��tP�d\��R��$���a��3�t�H�:�<�(��Xo�X�0&&��Ґ����l�ya�:��BT�I��5��EN)��J�C����� t�YC�����mAݶ|�k�Ԍ
.�4z�|�pM|)�L�Zo���o�v3������ˈ��ȹ� ���;�V�
w�,�]dը�EwK]+�d��>=k�
�>L���Ri&
�~X�R��;�	\Yn%XI�b��Ҩ��y|������ɖ�5�ٯܚ�T�	ǜp��G:��L*g�/p[�����E��O-]
nvqԬU���\�d!����|��� ��>�B�h��il�H�>?�Ⅿ6>�ݎ��ءqC.C��>�#�U ��H�J�B�#bB-�ز��N*["&z��(�9��$T`��M��o�ͅѭG�L�Ks4ᾛJP2�ԩ�����������(�40֓��P$ZS�^G�|rhmR���<���H2�K�2\b]nP��)ό ��5c��2׮E��Ϝas���j�w䄫S%g����;��`�&J>�'�	ޱ%?Z�Z7�� �3�r'�M�qH�%�����'	��D�����*[��DW��:����O�+���n��������tD�W��{&5\�
J��� +��^�)�׺�tc���&j���.��blDf�wѭ���r+e�`���}�{bs�
��I��㓇[�O�[K��] Q��~}Z��AG+,wx���u����!��DG1�-����j1����Ī[�i#��ij׿��5;��� �ӄT����w���K��*R�)�̣�1"���
xӛ±��,Z&���x"�Qv�,\�����!�$ٍ����<n�����[{����uN��ms�.f�bd`r7��b��%��Xe�1�ߩO6�A:_!���yw�)��X�L�f7N�G��b҈���{�)��Z��ӫc��fo&~
�[�N�`�x-��	"�����L-Ϲ�J,?��N�2du��$3}/����磷���h�0a��M��Oց��.�Z���j���2�;ۓ���ZP����>o@��_Z%�����?p�^���Ŋfϰ�Y�խ��Y���p������
)��V{)�f���ȯ)�Z��B3!\��4����x	����E�`��7��@��t�&��7	֏�ZޥO{TS�T����U
�B��*�m��=uL�~��rlm���_�Xn�>��[iL������9�W�P;����k�V;e˅:�ߐݲ�&���W8-$��B���R��r'L�˕�GN���2)Q�d����X���2�Ż�z$ �n)�w'�^�S���s<�#UC�sTmh�a�?m]�+Nʝ��=�Y�Zg"���6���#"pD?H��4�]<�(\(�0m����p@Bpp`��u������|Ђ�C9\lJ�?�E� ��Ҫ,W����v��F���Bj�4�_�������и��
�P硚�pRH�������a�����NO��doha�R5��nj���ag�z�Q�
J�(B��� b�H<{���ǳ�e�Q�5"��5�����������L�=	�`U�������W!}E�`h8�dS ��֗�����V��&�_C�Ƃ*f@?ϕm�5�w���w3�0��L��zA����Lh�RΕ`t1	�j�涀���s�����j��������� ��E���.�����] �-���s�^X!�+%�3H�8�A���������ӣ�8��L-?�6k��Z�pA[>�I�7�o�,y�^#7��5��e��������-���a~e�W�=R�j�4K`Vaoȋ@��V>��z��J����A�bDf��o�n�M���0�i��x��<��r�
)W.{��<�;�����Zb6V�x;���)e(8%XS�n9@,4��H����"��.�#�� ��c ��,����hЈ2�6,C��U��+���̸��M�1�5��CT�M�l��T���Yt�k�߂_���mi6�r��'��G��^��;HD�,��K��;FI4I��I�._�u��>& a���)�#Zg����թ�c�M����PP�>\Jy�:��묾�>k���:�PVs\�47Y�\u�au��M�?"ݫ�S������0�C��5!���ۃh�TPڛB���#�)j�e�PJNTud�e[��g31�7����l��Iyჼ!�6�� ���U��p'd�H(�#�i�ͥ����hs6fgD4���鯹���~6����c`�m�����Ȉdcq!���C�/f��[������S߾p�?��$���)�e��'4@>	�+$��A���V{���
䝦�:h>�B��u�hz�u.�eY���m2��I*Ƞ��=J͘ ��_�v�-	.in�k�U��#��t����y�P�瀞�E�v*JE�w�}�V'W��(�3�B���u��&�Ndԭ)���#Cz޶�/W��<k��O�{R�A�K�:�7L7*�YF���K�����6%��K��HWe1���؁ ��,��fІISU�W|�n���1��6qJs�ȅ~�l���b��!D��>�?�� \W�x��[�A)VM`7��?S|Mm@�޶hp���(-_N<Kb�$A��y�B�B�h�9�<L)�P�������9Vo�Jن�W��Ә#x�R��֬�WJag����g	b�*N�n*�+�35-ʢ�Az��>Xa��Hq�2D1�mP&�8�N;lk�D��2�%f�d�B�/R�}��e>N ��I��䉖kJ�*Zͼ����"
�IQnE��tMm~o^���5	0�iKv�$2Fw��kR�l��M���!p<��13��zO���sԯߠ0���\��$����~?5��W�zj�����>ԴT�C���l˰-��l�Ī��RQ�8�֐ �T�����Ͳ�3`x��,��Op��s�A�SI��4��R�*>�������0����_�&T(>6&��|�J��~�-��l'�pő�� �R���3�_j�x/ ��������SQ2�n�K5��굣�:�dQ�<n|>�����4��p�6%]u"y7n�=^:�&�71P��������W<�!�M&.�Ly�G�rD(Lg`:�1*�\�ƒ!l�var��a��&�g��J+O�<�\����)��t͉6��׫�p��0|�^���%����nc�#�\���K_���K��+ϓ��S#� �1�R�w����Z⨌��'�^��B�4"I|��e���[�$ʏT� ���T9��8�U��>�W'�w?28�D�Ep��.�c�A+b�ž�w�*�Ÿ�KK�|Q`'�ŝ��/�?�O���et��z=&�-�m]�͟E�R7:�������yl��5��īV��u��;�G�w�$�?�����R��OO��M���)�>���hd1�L�ؽN�����<B��-���a�V�gkҬ*��Jʃ�c�O�W9�Ĩ!H�>�Z��h<a�+ʿ+1��^�&�c�}�d�R­�nr� {k���=�g����r�W�������m�̀��r�

5s�k��3Im�Õ��G��DÕH~x���	��D���4��/��N:�y�_� �ƉE"`��ik%�[}��b�\t�0�:�a|Ωϩ[<Xoi����d���[���'`Y{���0�Q��Yx�g��[��
_�HƜ
���*w��K:G�Ȁ}���M&(�@���P6�M�� ^�IU�㭿f�
>)��]��L�s�`�I�m�\���4h�W�u�����6��,�W|��;��J����*�R�5������y\�pd���b�|~�n/Z+Ti^�ʹc�Tur��c��:@|��<��
�������dpcLԻT�N-�*ɾ������~����6<w��(Fd��,Q��Np�ә��8���Y�mi{OJ.�I%vh��?�t�5�Y͍���Ԛy}�F�b�b�j�5���6�0��5�e���n�M�p��U���n-IJ���{��K=4��/��l�msϜ�D_���Xաn3kga�H���-�~����߶�@�&w�%�\�J���_��/#�@ׁ�1[R[M{�RrT��}��E� g��Bn!"B=o�|K�b!�m���(�ݪ�P��-;wˤܾ �48G+����M&gos5��d��������K����MB��*�4AN�by�/Z#�]˾�o�-�@�g� �h4B�?1���B�L�б���`5�d{���D��.'��Z��6�
�Q%�QQ%���t�=J�f�p�p��_I�<����&S���g:*==Irb�<�D?5�Y��f�v�'P�7�>���܀Ӊ+O��,!BLhh��)~T���.K5�D#�/�Qͦ��{�}� @�s��h��&H�����ʥ�z���_�a�,�h��_>�l2��FD���;�������Q��>�q0J�W�O)�"h�]��k$I�L��[�+�T3�qF��� ��갱�ZM��R��l3�ۻɔ+��{E%bϚ�<�=_v��m��A�����@����/��2=��)ls���2�g�� �ޘ��+
���)}-h��ݝ �| �`y�)�ӑ��iz^�(�HPʢ��r�����CܼLIa)x�1�#8~�įV��L_�:V�eR,�g'�k�ˋ�_tl(�C�gQ`�(�-��{�	�&=�as���#_T�R�F�gCjA<7�nE��*P�g�o�b�pq=+����^�Mo����_++Z `�� F�Y�+|)ӱ��SĄ_lia�8�鶠��#�7?����-�n�����IÛs|��������٬��Q�ꤊ���4,�*�Q���E��pd�fQZ5�@��n�u��H�uN���:�;�-Ā�����NQ�
d����f��*�5��� #e��F֐Nu����u���bͤ��3��4Eq�{�_��브�����t9������^[��+O��<�g�+|��Ǖ�><�S����Q�]�f�3�`�T�K]y�A�K�v@+��������.6�D���-4�b�����z����M�^��6
>pm�ZfA�NM��s�1����-WG�)�[��C	l0"���:�T'Ie�Ry��*B{�'_��U|�Xio����a�_�t;b���v�\?�_�������ƳZ�ӕ(f�N�p���ة���f�h�0��@�q�؎�͛a��Pc�ǘ�l2�[+�=S�u�~ �E�B������㩭r`�-�&<8����(��̩X|H��	p��i[a���Z��&#���SpL���X�ҏ�
\�SD�-YJ6�!Mj&����f�f�bH�����ӏC���ሙ�rf�� Pq���P��"f�Ϙ����ڨ�L�SE��N<�O��1\v�si�ʂD(k���t���J)o�}���e������Jտ����C��"@@x��[�eM���4�r��x������FC/�޷'�j}ۧ��DaeE8�=1|��k���r4>H�@��6�j��Z���|k�tΨ���T��Q�v%�S��]H�V�~'�X���q���n�І�0�
e/�8�m>�������|fb�s'��o�J���]�4�D��(�%&؎&� ��MʮX����X�úVwz���� �rA��>�"ݢ�ª�j��dDK[p�`��fvu(���0�1���p���]בԸ�����h����ݘ߇S5�n��Q�)��#p��2ْ!ch=�"�7HA4
�W9���8방v@���2]��[� ��2&��P+UR�# �m���J��-𤓛C'O�ǚ�g��cxV�#1�>���H����d{㉡U��֑,$6����Q�|)���ᖏʾ5M`F�.HR!��k�Z.Bt%O'��l���Iȗ~�1�Н�C~��v�^�dBF�1Z�LTIs���'���.��/u��-��mY9p���n�~D��>Zr�{մ��ˢ<�	��̈́٪X�wm��<y���?HE-��"�u�W��0�-M������ŀR�I+�����~�s�bG��3d_/�Y!G����*Mʯ[�O�?�������-�dD���qd�^~�_,M~ZA�%����V&��ְ\�}�����l���Z�qa��.�ע��|�rd�>f؜$��O@�܌E�J1�>���G=X����yu5F17%B C��BX�>���o:��X����i��BC�ૠg�/T:t�p��w,�{!���q{.u�5N�"?�8���V���d0��]�|��jRf+�¯H/�+�7Q���A�x���2��!�!�s����bg_8��3.s��I:V��oA-�a���&9iQ��x�����2�*�C��`D�e&���G��f�2��qBo�T������g��N�\e�p�~�	�L������M�AlR�1��<~U��pi��B+�i<������<�J��8ԅc��CHTu�M[I�,{��ZO�w����O�8�һ����_�
C�gpD>��Tk��b홻���p���X6�&�G�׊�$�`=2��vƓ���Ihs~�:�g]c��L��cO$���G
�zA>d�R�~������R��ؽ�Z�E��K& ��tp�~���&5bY��͎����z^@@7���V��꒚wt�~�Ro���z0�n�X#�^ŉ����	tx)����͜69x�I�q�t6 � ��(ރ��g�P�%�a7Ă>_��~+���\�+�&,m=4�[�b���-��H@�c��֭��ڃ���<��m�%�1~�ZS��'�|P�#��^Er~t��	�q?��=��M��.L��P`�2��dt&��,(��s�t7}�g���X����αU-�T����R1�V����u������ϊ):g������[>����P���_���ma�S~L���c2��i@�i4� �cK�q����Յ>�O�p�IV|�v�������)»��*��B頧n�hG>�{|!>b�����TčiM����ϒ�Y�!gL���D@���W���w���5rN0 �i��˙�(�q�R1o";4_�>��7�#X9��{w�
�����?���!I�$8�b?�1}5ê�Ƣ�C����(�Si����D%�WsU��<5i�d ��6E��P�4���\)����� R���Ni]Ҹ̛�[�Zv�-<�������D>��)�ù����h4b�~{_�;*�϶�)C�>���|�U-R�+��l[�9����je�3.�Z��@��>��5��ws���l�!Ȅ%�+��Y:Q��?%z-|�)E�H�4u��y�/�?:��A�W���J�xk)��ʪ�7q�����m�o�P[�MYwsR��U5���**�As�fP7�b��8#5L t?��@���hjL�f��́��4�}�	CS{�0�澑����wN��_[�*>/�dOS�I�G8}�ۮ��(���.~����ai!`��j�V�@;3��4�⁴!��d)�c��z�����ľrE䙡f��79�UQ��9��WA�z�A�m@3��)KJ�n;A���
ʒ�,/���;VԲ�@���`$'���4z���QQ�c�~i8զP���Y�w.G煩��i!O�xE��-�A���l�ҭ���&3um�Jx��pnD��&�Lk�Y��Z:���n��J�}�^�Y{@�nƤݽ�ư�C��GZ�����x��
��'��a���-/Q��j�m�,J��>��3~{�H�q��(~>�.<Ň	����0���Yԏ�(o�R�X���|��!t�2�48���#Dv�\�Z����h���A��E�J�3�G�������0RE��y_��Ϝ����5�7���jK����s�ׂu���K����|o�9>�P���X�BY}��9Au؃)�ؤ]�_dC��sd�/�z%~�-�ta��i���T��Hb�j'3�|��E�7N:�U�+�,�9�����&�K����6�Lc��c�e &���?�˝���< ��eK��L+	�}�0�i�b�F��&7��y�[Ǟ��$����!x;P\~�Nq>�;�)�p\d\�$�j�7r;�N@�:D93���~nR�����Κ�(�4���3�lH�Ӏ	w�`n��/��)֦�v�y�WI��8h3T��D|��8�0�_�k8�`��qe�~-���r���.��p�J�A�V?���gr�fC^���ɴj@���V�2�CPI�{��i����mt)Zf4�F�v�P9C�jI�A�($��@	�V$��TB���
_e�2�/0j���&���@��vc�z�+����6���?��B^��r�8��b����ˬر�{�B�
�"(�]�9U��v�X0�<s��`�Heu<��0�SR]&	f�ӱh�Z�*���e��9j<&�h��bd� 5��A���{��Ge���d8�dn�2�*I�x8Hp¬��}7^)��Z���څ^�j:���e�y�N�$��RF;u8�l���WJ�-���������D�����`NOM�l����ȏ$��A#�D޸���闺jr��.����(��7�)�Ċ��~�0M����ҋ���=oXy�h�w��Vxytӫ�3�k�k�O���4��3�r���f�=��eN�������XX(*�g�E�k�T�,�~6R#�gb���,�aCc
2��NͼN��d�\�m��+(ej0��k%���q��X
իK��N��s�h&�6�ؽ����`5ᵦ�lʪӥW�*7��qf���������T�G�0�{���ߊ]
N��M�;k�:j2�t��h�g�zk�dӣ�}��p^���� �:S�	�a -��6�c��G�`�_�is�<m��?���6k�yD�-x+�QD&�i ɇvXw�aU��ŕ�2��#�^�d�s5���K8C2������)\��K�ǐ�N@	��۱2ջ�X��EP� �bB�|��S�lX'���}?߸�u6@�0j�S���2R�V���ŌAR6a/��zc/ �k�D����u��6��0l+'[̺���9j]�=ӗ��M�c�{玂�r ��B��H�@QU��H5�*![E������(�����4���
)���Y�N��u�I�G��X4N�9b޹��Ϻ����V+�b�<�K`��A 7�p=0L0C	�2����)�J���y:�t�͠U�ܗ����`��PQ ś��G�f��~|z�؁�6��$W�4�r�s%�0��-�i�]�x�V��}��@�� ��
�����Kv��Ņ|lo�u��*@ZM*(�%�C���^��Uγ�WO�U�7S���X8��4c�_ s�'�"rj�Ut���M�{�t���/��s�	Uf%����+�E)|�����Qص���zZ�?Թ���Ɣ��[\�,n�a	{�Y�@���p�8� t��{���"��6S[��3�LP	bI�.�HH��,��f�q�DF�E���	~8�hW�L0�Iz��ݝ�~��[��_3��^M��4�p�3�! ����I����㉐�SK�J*��ŁE$�(}�>z�ĺnI����}�~ؚkn�����}�W^T��f�
R��ML�
z#r<:�T�>�5~�?Xؼ
�9���Cބ!P{�!M���O �����b;��)�J{��<��q&�+�F��ߩ�k���,@��� tڀ�ΟK��������y=Z���@'=�9�辭^��@1&J35�ڇ϶��d����KxA���S����_^L��	�=C L4��b2�[�F�T5*���4�>u���8U�~�k�jR�\�����]lJݚ0�6��� %��?�����<�ךb�y���&:!ɸ��g�4 �ljЭ�ZV|���6�͂��2
�$�S� x�oY� U��~�?ā��N�>���3/��m�g��jn�1B��u�?�!��!����ͅ��L��Vgڐ9'Z�{��up�'� ��������2�~$��ڔ��`��G��[)Q}TB�c1���qS6d�͇��XL;�XWf:4�vHt�~,S] �IDBٙw�������K?��Phz�6M��ed�
!�Pa`H�L $~�l���)����Q3������VH�ʀ��A뚩�C�k�q���5.�A���:�'��[uD�'>���i��嶊��8A	ZD��1��)�Y�g�_1�=���:�lc\-�!�����u8�+��$v�ݻw�ԃ;�VP���PMhE�Z���㦺�aG*!�z�z���m�g���ǚt����"q������[4. �؋u���[!���Y�����Qc�>�mݴG�+5c�P'�E	d�`�ɘ!�͆@o��B����q�����B�<��~�ō���3~DF���5}���q�L����CA6��ս��fD�,�{r��Z��p�h#��^+p G���@䐐��Ֆj�QR+���5���g�"��2���w��9����?�����8�U�V߹�b��ԛ��������'㾐.<�%G��~���rq��6y2G��eV:9�@� �M+4:�I��D�bY���ȇ�J\�l����Dw@����l��#my�p=J�A8be�q����P	�A��,���xt����mL�';�H�+����]�j=�#�&�������w����R�\w��&ln#:�o��U2���)q�gX(�.�l������Y���x��(����0�bY��t��˲ХD)�k�E�����=�d�T�g�wc��*rh�h�wq��ټ��4�*�^Ha(`n��H�_L�Z�-��������i��K��8������3���J��!�F�]N7�rQ6>�d~ ��7;3��c��c#���� ��A���b��C�^x֠,=K�����>祠�o�¯u��e��@˭��V�<3{��5ʶ�y�u�F��9.�4���ɺ�����fp�&s�E��KӺ���\9��@[�O;7�x�����<�;�<��� ����.�wk���')k.ά����M#P|p��,x��b�:<�����h�$ߜ�S��0y��G��$�Z��4H��g=h��1)K����X"��/��{P(����Ş֧�o���/{j�i��*v<��:�h�Ġ�e|g��%W��17�y��(�8�4�z�J���_B�
mw�k�n�h�]ymv�@���-�C�7�{�ŻM��*By��
*�������-k��f�S��>��L��j��[R<�+ x�y1�_����XG�GZݲ��r�(����>y�[��-\�sЉ�C��¶�R>#�����/�fִ� A�J֩�	�V���揯�Bb���o�؀�h�~�G�(fTA��2\T�q�?�;W��>�	��b�Z��D�g���^nhy�b�ݣ�Dfi��E�ƘW$�-�8Df�������=��Â��^#>�$S�R3\7��zyě��M�	،z^���.\�x��T��D��iH��`�a���l�wk���ӈr�o�&��4N�P�Qy�6j/7��K|	�w�8��T��c�)�ә��ց����ݬ0tœqU@��4�D
c����@X�N����?lT�Y8_�yr-znr������Ś[�0��Z �&<��"x�T�����S	��{��}��x�MO���2�2z��̲T�4p�M2)�� UZ7 1�N�	�� ���VOr=���i���
x�'�}g�))�Gm<�&����n��}8��R�W�xO�1��L�߮Ux<A���]��\��v.Ǔ+� ���X���k����Y,�?uꆼ�u"���ei�Y�"q�l� ��V;�G�ͷP�h'�t�R�<��E�#�ȕ�_�v��W�4�d�S�F��pdE�y�̜����l�%��_��>[.��ph��D����Ds�mC��	�t���bq���Y� �����q���\I�L|!W2w��Å��͖�z���'{�ՂAT���������D�M�H����]�D%Q(��ˀ������,X<@�V��FW��b*]<�n��O�����8jQ���9u0|�����(V�d�r�z��4�'�����),"�}9�CC�����v[8.�ҖĖ;8�T������d��Z��"����H��l��=�?�M>c��X*���t�-����?m���Ѱ��z��cm �x�ε`,�/�<w��4��3��Pٲ+�v�#�T7�{g�-�@�f��>���PЈj"����@���ڿ�I���?dG�#�^�LSj6��Z�q�(�i�j�p������k�;�Z�5m0�T��V�h���j@�o�٠ݣ�A��Ua��ۍ���ל�C�����ѥ���2yc����7%~�*"�����Cv�)��Fbl�%Kowr/#�Q6f�j�������E��--V�x7��>�ެ��T,��}Md��:�.���L{��߫�]�{ܨ���K�L���� f㢵�+�
@�m,-�*@�/��U�[��Fy��ڲ���0(����4�3��A<3N�~?dc)��Dh\l(f�����֌�>�����%����D��*�)V� �z�%B�̍N&@P*0���#�s#xQ��z/J1���Y���yHXc���7�a���a=<=�h��0d��E�<+0h�6#�
�C|��D�˴p#�5����t�Z�X�����8�D/����r�4./	�_XX�R*���Xt�DV����b�`��5W`�}{*L7V6��`-�� L�UY�T�Y�X���+�C%:�� HMo�����`Ψ1F*��P�F �-޹�������O�@�	�.[�a�,���K�S�kƱ�)��j�qڃ�೜���^f�m�^�ߒ�p
Е�o�T�t4nP�j�q�K�@�9Ǭ��L��.7)��FV��T�čc��l>.(������V�ר�S��p�
>��з�:���}�}�3ϐ�_�-�p�`��!��v�#*ĵ�9>O�	���}E3{&��>yd|i� ��ʂ�^�ż��|匢��E�:*�j�4��&�~b�Z��+�0��Wb`����S0G���J(��3pMWoq�߲��U~�'�Đ�Xf��|���S=���P4C���խ�i�v���ވ��O6]G�b_n�Hk��0`p��NH�]n��,�u�˷%h�z
H	��%2K��L0<(��W�,U��qI.N�2���j�N1�q����+<<'4X-�+�,vՍu�o�+\�6�W�[�z��Ai�� ���/�:K�5�N������J������K4v�`�ة�rz���}��`ȇ��w8S��-hS���oP���PUOʛ�fXɳ��7�a�U*��4e ������b7� ��j#��'�Vzb���ϑ]k-����u���#�q�~.vD�ԍ:�Hh�6�w8��a���f!��<��*���z��_�~��&*��!�L53��kb�i��.�������9ha,�LH�9.��̜�+���Ӭ�0�B<�����\�-���ؘ�M�Ipf_L�i�M;�g}!��hɆ]kF�'ϔ��!Jy�%	s�M�T�3u2��ѨI��YJ?����}���ݶ�h�4L.��YE}��Q�������n: �(�?�)̺��劊�iP�����(4�Fp�d�1g������+���57�	.�F��PX��{��J�|(3xP��~7��`�fy؍����� ����R�1���#3DF��~mG�=/��J���)�W��p����P2��D#GG��=vR}ɾ�6��������+���,}���Y���j���)j�[Em�1���|�I�(\54�����d	�<�"c��vC\a�>b�i�t��t���%��wW-;��rr � �����^R�CUT�r���[����lQ��K�rI?�InM[I����x�׃i�$�qg��(/[c���yt�_6k�?t�1�i�� �_5R��8`��R᎒d����x�y�����Ǫ�(r���vZ���.a�w��CLϷP�L�Y�u�%����OĪv�\�CП�U��DA�We �"l�p?

K�TEI���v�b��۔l"���"dc	����*�`"��։��`f��f]i��Fj���<G���%�# 0_3J���=έ Ʉ7��Jֹ��ǒ'1�n(ЎEc\���7"��CM$���5��[1�Z�0�R��+���8k���I�W�F�SP�#r7�G��(�W^1`<p��g���������Ԡ`�>��a���>�V��c�vJ�
V�cV䑏H���]h�ъ"8��w5g��m�h6*�K�BA_g��8g{���=����-���wւ�f�=_{g;(E�?/<&a2�f&�if���V�_:�
�!T��u3�-`��W"��탔A4h�j����jpg#] �<���4�W[XH���?�g\2� ,���GS��@<� ��l� �|K� ��kCթp�]x�N��g�(�j��p�;�q�3,bֺc`ZC! i���a�e�� j��g�먖��w*���\�,��$.���Nb��(�����_#�l�c���Ɓ�d�RI��Yˏ�R����ڬ�bΜl����j�]�i�QO�+����e�V�����&��c�;��,�,v���Ɗ�]��	��B�*�@��bJ}U�T���N��to���|���?X�:���٨�f�v�Y�E�%���$Op�XD�f;F��wq"�Z.��
)�F�� &F�dܢ��m,��"UD�� ��{RXQ;����r��_�[��b���[��a���`T�:IՏPN���p�T���7�я\�=n�]-��^G��|��ڷ�h���_��?Y�3%Ȑ��	K�l]\�p���sr,���LM�8Јhb���Ń3F�bF�(?Hl���F�ڃ\S{w�y� ��`V����j�|.x�<��CS8���zᮨ�4�� ��y��8��L�-��(�|1��K�c(ˈMɿ*̌4�����<&�Z?r�w�pM��Ut�.4��yb'�ZR+3���������|ÒP'�.��Ԗ�"�?�5q��gQ��z"������dk�^�n�|�k�1Ј4]��!S��p ����ԈE�?3Eǻ fA��#��h��a�*[y������*%����е���4��u��$"���2n�^�߿V9�Hg�g�f����k#��_	����S�̞s��?g�������$TJyπ"'�dEm&�������3���e�N��[�b&��=:�������8���(��y��ɟ�|��?��G��\Z� F&`U������.�^��������r��:د��[���ʱ�Hs�8���e��=M��F��֟[�Li}=Ĺlo�~Ti�)�~��,���kr7L�7%��/�p_�N�wN7��2k��C�,F'���ɡ�
Nq��LW;����@U{4���3���8�Ԡ�ȟZ*o��ؔZ͗�>�L
� ZˉA��	��G�\\-TL�ϕg�.`�L��R0��ª��9+U!Z(���ڏ2\�BƦ[�u�0��@�v� |���#p���u4O��:��(+�Q[h<�kz�9��A0n}�wx
#z#�:kz׺����kyO���iV��<*��&p��?:��z��/��R,D�Ua���ޝRQ��`��>T�dlJ�A|]�E��֯��#�	B�E בO�!���3d����`a98��0m���X=/��ٻ屜�ާ���7�-�	d��T�Y^�s��5c�)�"k�&F�a���ލJ:�ed?e��R�BM p�q;��o?�7���<�������bʓckNگ����
��!o��=������L�Cy��T��{~�N����[i\��K��_���_�$�D(l�ϩ�\�	����*�/pg7,*Й���T�X�Y����@Ӝ�;�.G��_����mɷ�.��!�gby���eV��ٗP��u��*�s���/��t�xY��\5��LR�]��kh�0�\�����<��X��j�xN<��a:%c�Ub�h�SD�nꏅ���'�h�{>WVAI���_��qQz�$���%��0�h��<(�:1�6��~��ޤ�|:9�4�K��B@bsɷόĢ�޽�,*7-,=(Rz����=G�oҮi,��3��,y��U���MMl�Y�Ӫ�_g,��$���~�2NSx���cY>�Y��U>T��Zr��y;���k���&i��=��(���{�1z�� Wc"%]�P�W��d�4C��|qi��'.���VP �hC��ZӱF
��l����-�m��Z�?8	\����wM�JÖRXf��W��73��G�B^vo߉
�[^��h���D�����|��Yv�D���G�tZ�d��ݽ�+���W�;N��''��EA�U]�7�� N���&�׼�7j�Z���sp���hQ�/�I�Mb���v��}g��[��oV�D�KK!>��) Ǽb[2 ��E�+�G�Ȕ���s�'RW��X�*Үf�"�#��<�s�ýʾ�qȳ>���O@m���ix�:W�]�tSgŰI[�Ϊ:S���Z8�!{a=V���U��L��۸�����I�ܥ+T��&��)ߠ%1��Gɕ!b�&6%~�>`R���~#�m�yR��3?�x���g�Rnɥ�4eI�������)PA�����F/�t�p����[y#.!ʁXG��i��}��\=�|9%�3�����K|1G;s���b=��Y������^�7��$�oBc@���0&��99|`�1��!�lv�L���R\�����.���,钑��l���u���~�]xB�~у�Q�v���O�;�Ȉ2�͵	���;�K�<�UՀ�D��6-�������y(j �0�&�C��9"���x�E#��a|ۦ]��1��E��M�RcvHI {����Y��5D�Pw6.��Ư]���oSiJ�A_�\F�����m��8�Ijj�n�n@~�QU�:�H`���⌮+�,�7bu�t?z
��^�(��}h$3�q����}���i�(��yJ�*S�o_v�z՚1֜�y��մ=�xYD�E�.�-�g�q�E}���nI�	��=w��P��wl�r���R��O
D��5y����t�Y��"�H +<�u7�|�����qc ��������:�{��cs�^u���=�lE�N@�H֤�Kk'A�r~�j��Ϻ��8r��Ǒrh�y<$��MW���ld�B�Iq��l\���>Q`��s]b.�B>�hu�腜h�@*C�%#�Z"��{_�s�G��x����:�>B.Q�-g򣓧�_��SXTb�}o�'�>��,�~���WMRa�Q�h�=����,CX=��<����ݐ�852��g�vB���Өj�j�\�M���ʏ v���3=H�4��+��Jt�P��w��D	�K~�ј�C��/B6@��X�_�A����@���1����:�Pk:E{F:|.e�!5�R�B-��$�]�0t���:��7��[���dvl�R�jhl�4Og	�.��)b�!�1�m��
W��- �b\@�r�`���yLۍ@2�p�#������Z*h''Z!W]e�K	1���o���2	d�W�ҊsZ/�\��D\��?w�%�ԧB��%��9�	)�!æ�ް,p�~J :@I�i��Z6�6(��x~�B�ؗI̫{��7�cC����|	[��G��0���{��V�5�����YJ�Ā�R����|@fȃ£� �<���u�H��+|C'�H�_�.�c�I#���,}\��S��0���+�đ����;ٝCl�02n|���K:u��]ݐa9��E�ħh��X�f�%[3[���d<EB��|��%}�E�E�)� �W�*�.��?''2E��`����.�q�a�IF�v��q\0���H���t�u�"��0��G���'8?�����]�+/�
S��M����Y�
{�oC�ˌ� /Vz��ez�Md6<e?�W����fA�1�x������P=�)8�B�S�kSK`##gwF�6���)��֨v�b����8y����	E�ڜ'��g6p �o.9��w���;����:Ρ>���G#{Q�|���U�I�5eLNȺjz��cbIn������%;��������)GE.g�~����W�O�{!�>5Y�Tev�ӆ[`:���%g	�G=�W��cJ ja4��p�6��Я�;܏;. I|9E7��0��������t�;�N+qJ�JS�Q�� X/�Ƣ��,��v�,J�y��V�PW2o/)N3��wͼ!ڵݚ R��q*"B�g�Hf�Q����h�4�[+-ܴ�_BF����4AÜ>iM�O>�(\61��!������-Hjڂ:c� Jm<�RW��z�d���k<b��IJ��O}E�d-�X��$� ���mU2:���[�#:�"0�_ϓ�@_j��AD��e�|2.��QlD�����^\ ?��S��{�*Φ��x6X�~+�o�MF��)x�U�~��_�$T��J,U\�R,>��<��h����[�E0��-�Z�����p��lu�zm���+ �P4K�
]vo��[�U���ە��LRcjh�c������||ȭ��~O����@+����)�	�=c�;�Z�_��*�B�ǒψ#1�[�R�?r]��ScgChxI��R�W`,фJ�����Y�����~�<b^��F!��'�[Y�#��op����N�B�����O�ʅ>���+i����B-�sd=sz��o�hQE�
�\E�}�")0T�r��6Ӎ?)�'q\�]�)�3��g��~o�;t��שgQ=e9#���@������Ǎ�~=y�������{Z�
��f�ǔ\�.��^���$T���_9�V�q�?蜈�j�mD�T'�R�
��N�%�<1�͚�F،"s������i���Y�0l���Sxur��qs�ywQ�YeyS��QM o�9ϓ�d>�_m9.RfY���� ��C)X19ȩQ�V��dD���Ŗ�U�z�K���'p��IJ�:ƴG֭t�6aC�]�J���3�$K�>y+�{� Tz�Y��N�*%"� �3;����`�{n���J����;���Fse�9d�ǝ<�����g	��`b:C�4F�c��(�����|i1(2�Uwl�������T䛲"(|q�煫�j���IE�hʕD,�3��i�lpMc��́R�	>H�Y9tR�X|�Sl+3u��@PA���gu)���,!ő`V�\�<�~��t��:�B����M�V��'}���$����_�P��K�@X��l��xv���Ʌȡ��6��ls�S�Ny*5|�Hγcg����@���ԋ��T��c�����)��a=�����+(~���+����-49H���+�{��;�f�C��N�l6$�nn���F� �`R2V`��P�ֆ�O��� !@~d���*�=�� �-0t�}��bH���������Zo�9>��)�z��s���o�k��8������º[�T�-�KƬZ$���j��!嵒�f�*y\�x(<#����)�1g
}6�0��9h]�B寂�-5���'E1-~(�>�l�z�3�,�}K���;�� �.�O��*�W���b8'S��FO]���K��o:G:�f�4����U�
�CVy�&&9�!��GT�_�|1�����#3�����{���WLg`h��L��m�G�v.���������l�q�P�|��T���dL���֧Y\<�R�)�4�	!��_�����M�.<*}v"��1����.>ڄl��|qTA&_��T��NU�`�5/��/�b�N0��+�3,y^uI����ðN�r�8�s�HG��L-�3dW���� �^1xnFP8��Ʋ"bn7�y�������s(7��uTV�Oe�`+(}�XKI�Y�R�qñ���?o��F"��jp�5�
7 yRf�R�\�o��Z��Z�Y-\|f�}#�`�6�_��{� ؝��F׹�Bx~g\��$(#@�q�f��g��4�sr�(�_���rk�ȁ����(�t(����W�ś�t�q�����F�1���P��[���~����fO�gY���y�+HVdլ�g����{�B��F�E�Z+4g�=���B�5���=R�L-Í�+�6:Vn���:l�����%��6Q*t[B��հq�9�B�Z��I��������O��vI�{�fӂ�ΐ�=����ZG�_>�m�����$�Id.c��E��)d�L���+ٳ+疜9J���'��;ߑ�(��]�r���o���q^��(_8�ݼ��:2a���z�*)��%+�m6|��ܺ��lg&��� ^8s���\��c��H��T�n!���{�E��ǩf��`�����l
����2���ς^��J�o!�Clڢ��<5SZ/��͒�������F�~��2O�(5�Ep���-���c��H ���E��+��,��]���D�.�;��*��Nx�yNS���e�`Z�R��]�T1��C�u�5��k�_��w��ˬ��8t}��r�x�ݱnw&v��K��7���E{D?!�1�٦=pj<*�e�D��˿BMw ����O@HR7D�n��b[�E�lH�*����g���'.e�[�z�s��XUBA�������C�V���H�'��;�M�z:�9mm�2M�{��F��B��+Y�K���O2N*a5/$_��p�tv�	Gn�Qq�*d�>-�n(U�����V����H@��J@)��@�ʹ�9g�O\4/4�]rn���:����U��|6��gQ�"��>j�ᆇ1�|R)v���Bɵ�ʇ��e&(�>���yd��#N^_s� �N,�����5�\$�m�����&�� ����欎REhO竴�r�K�'�J)u~xa�y^����})I��������_�,e�%˿V;�00s`������y���<mk�� �z3�I�,�.��?9]�/U!�7�m����/�k�05T�4ʀ��\8��:ȬC�Wz��ּGo��u�X��BHxԗ�<(&���>�f��e�d�H�|l��r��/�A]ӽ\�[S��m��L�"	nk~.>/��Vhn�:���('�r�8�� ����ß.*PjWpэ	�b��f����Y��(jb6,��щ�#�Iѷ�'�&_/������t~�{�?���js^���IOS[wKū�<��5~b�J��"j�BD���2ܲ_�����r�7E�!c6u������q.����zv�Y kAH���.�d����:j�(��o�B	�}T(�޺�<��(_�, �VH�䪴�x �a6SNAɒ���5�P��vsZ"_,5�k��)�z�
���������۽VW����|���g)A������s�sc������2e=��ja����s�R�sT���W�_�ɻZ���Kru%�t�]�*Q�˼�D��pi��B�{`XxE�Z��L��*�׫���w�p�0/�z�4��&���Y�c�en;�����X�W�$=�}FB,�	�x��v{�{� ��	��K͚�SHLr�����(��W�x��݂҄ ��N����ZA񩻉������߰��Uu��p�#��T��%!Sl�Ԗƫ����g��O����`�d 	��6W�?�r��dE<��[֒�KY�ȑ�I��rK��$>�Z%�6'O�/AT���}�}����dp���GV]ɞ���x�#1�s����K��n�s�} �bJ�WF1:%��]��|���S�Ϭ��|��CZ��tU�;-A�ܺf���wzid�l&�y��S|�(�%Hhd?G4u͡܏/DJ�G���1UH��I�+ס�oWC�\�boTzى�]����2�q�l��w$:��;R��J'��[��\XqM -��g?o-k��-�)���[�R�����!Fve�BJ�D��껄i8p�Uv����s��+_��x̳���gUOr�X�\
	_�1��K���M�@$��+�ԃ83x�GlU���Ni��1�@�����"p�b}͵�^�1���Z��E�~4^HE�^PA9s����]ͣ����`M�@N�����J�֡�AW��Fz���e�xR�O_:��[��3^G����������}.�Q���
�?A$�QIf���&�Y/�����#�n��=�0��_��$YR�g�&���5�ԝ�]m�q�:I(Ӓ����f:k�u�,4�M�Ǳ
l��%2�����D��s� ��:�܂?)#�kS��^R_�0CqOҺ�U����x�;��vj2R�$��8C�m9KA}��Q9pV���������l���r�F��MG��[vZ�*	� p�ٵ;��K[���n��v�Sb���x�։�p���=��e6�0���)Mf���e��ݚ��J=p_��_: ?%g,n�c�y��e/W,;'Q�)�8�ȉ"8C�e>Ha���u$�m;�!4R��`#O7���eB4E��m�wﵙS ��|��G֌�M����bM.*ij(�x4�w���)���F�s���Ys�|�?�}�C$0����M�n��b�;��ڪv"�g��d3���h���]@)P�#��6�����>�����'?�f��,��ݙ0(�`9�i$fUbF8|���{��x3m&/� .����Mo�Y?���}�=�.���(��	b�d�X����2����}_�Y�fب����!��ϔ��zZ5M� �1F~��A1�;��$�A�(D�g(��]ZޱL��ƳCQ�̱T�h.�kYӽ��<�ܱ-�NH���ζq����iHx�cb�:j��3mN���({E������%�y\ewL��r�>��*���\�w!ʽ�˺jᏊ��ƹ�l�&2��
u#ò��dw�H��� ��X LtZ�����WL���Y�&���JG�n�pj��_�{j{n|��F�*��Y��@��J`7�h�m�41��9�,|�6�כ3DڝM�����n=�ݘ����� e�L�(*I�k���f�[���}�`�5(���Fǻ�0,��O�}�{ռ��&Ry %N�-��,o�5����캎��&̔��K:��("�O'�����҃��d^�N��A�5���{�c�e��fiDaۨFyC -�C1�d�p�b���yQ4,V�s�K�!D���Ehu��d�j@e��#'�y���*UR���N����%̯΅I�������`��"�g��wq*{�L��<�v�
�.��1�Iv'�
.< �=�3��7�:8I�Õ]g�B���t0��o}M��#�mA	��v�\Q��C1ՇӔ��2ܘI�������LC�S��R{G*�ف��`1��m�2X�U��q\8l�.OWlNQ�Fjْ�H��G�RR�ơ6r�Z�C�����U��u���o�^{+�~_P@�������K��,��w("?�,��<�d���D,�t�<)w���ڤ/�2�p'Y�;�?^�xb_4�\:?�8�	�3�X@������oE�����;;�O^E����O�7�Ö��9�o�@;N�d�'�`���J"���=x����p�xb��r���E�G� � T6������;r^�]��f�%����!�D����e�KM�F�\��EXc�w{�[�g���}�g�[��)��vk���Ο4��]$u���
m6���.Pф����\@�~;���O?7�� \[)���:���B"��fqJ��=̋<0ꄪ��8_3�~�uRe~O�����P�Jʯ[��0�a1��d�o��oNvх��ג:4p��Z�r��dU�5�n�	�J����r?���ר�;x�oӈ��nb"8�|_V��J�ܟ=_��#��	@�'�g��H;e�H�ӿ��L�Jw���M�Rw
���_�iF��]��Y���i�w�U�\��[��˙�ڻg�� df�x�ƛ��I�����b�	+�O��A]l� ڂF���&̕���)�j_NP�|����a�Z�9�v���q��/ϝx���\�
��$쭢�W��sz�]�
�e?G#����6�U:cK%0����c���ج�L�Pw�(���K����CU�h��������0�Sͪ�:䍭g~�l��$p�E���7X��.�s~o��;��kz�"qq:Q\���q/��Q��$a��Wz�@ �x����e���Rr����u�t��l��Hr5�b1i�KCюD27��v��D�x04���[� �%*q֤\��wiJ�vY����#J��_q��ܨ�<F��0�����"���_����T��+p��ҹ��c��vs�&����ZB�T�Ϧ��tȦ�%�:�LD�`���P��!��_����g�ysP?\H! i���O��=��7�@"}�g���(���kq*M���E�"? GE8a�)����ͯ�4O�W�Z@�_�ֻ�m�ڊrL�N����&W��)X��NG�4D�Sp��Ű"��pLo��|���*��8�5f�4������Hx�*�d�g3d{�����so�/�I=R{Ho_!��i�Y	`;N1[�'<�8zR�9aiZ2���H{R	�~5�[����=��@��Ά���sȯ�(�Ii�c|~p+0�Ca��m�s�G!��5	��F{Є6��ƀ��Ѐ��Fe�^$���'� �z=���P��ߛ���1>��Z�$(�-��k��gp����#�ww*V9.mS�5�tͱ�T@ʆ�m���3���;��N� XbHP�ثM�ޠ���&	(�v
�q~�}�u3�3޶���b�CX�W�"�z(�(���qˁ���7��[����ܵ�g}��P_$w�iXxԹ���1��?	��Q��"u�%�؟�����+L:��+"W��5�Fl�?[��,aX���A���$��B�����\?�� ����K
3��7��̷6+;7��A��:�	ʦE0�@�\�U �{������my� ��L���u�xk�JQ�gg�l{�,���	�m�	��(���|5���)*q(�7�k����h�S�D�j�,�p]��pίq���1&&|���`r�5Y��Q���+I���V��A#���-5�-���F�{��/(���jtѤ�n=8����J��o��=��Q���v�Z5����@]�S���F���k���R�T�V�ja�m3��C��L���ҟ�GC��YBHT[���h�;�.��~*�p������� �\v�	Z�˭��?����6��R�7�[JY ����R�$�R��L�ٱ�6`�H�F2��H���h���+g*�_��2N�����A��+=�A*��xTM/ȼh�%�(슏�0��O��ϢSf�A��tq,tu����z&]A�%x��=�z�O��w{]���n�w����<�l6g�̧7���?�jN4)L�*Zv<Q��2�c�.1Kb�%a(/X�z1�ʘ�X8����M���,o%���X-��[��u����w�v�����1!r�����L�ilqFY����c�:p�̥��΢S1ѯ�Dx��'YnD�Lߗ��L��d��-G퉈I�t�?�b]�0������M�C��5����Q��� X��2&��:M�D.����n���!�y���r�w��b1nQU�W��	��u�<��0(��DO�1�8A�Qz(X����Q�d	H��4�v�{N����k�o�r�R��_rB:�~{���������p���~��-L�x��I)��kY�~]v����2
�Ac�0��#�
M-1�f�?����R�y'��y� 7(AEnm0��
��:�@�OţNom7��9O���9i@3qr�����/^�z3}��65���>�2{���"O.b��I�u�PBw���6hP����P���<�4~��������+*���i7�D�n�]o;>Oωg4T�}�S��\���;[I�K��u��Z���x޿y�&���9�����4��3�:���E֐br�w�N�[l�c�����g�,������J�J,�N����#J�߱�:B���Vr������^��@x���X&��y)��2���Kt������3`-��hnw�7��o�Mb����!����^�j�6Uo:5�rM۹�dC^����y��J{�zb�������D�7�[��h���J�-�yģ4������ �a��7��P��*R֐�@� �p~1�_�}�,mw��$�S���@(ռ���)H��T<C�\���J�f�SS��7�3T�)U���Եd+u��ڷ�r(�Iqk]��O�r������W��S�%oxVU{��ķl�0~`ʹ`/Z�6=���ʡ.U�g���q!�`3�w��[w� zp뢭pm<��!5�U���u�V�[�G����b%�@kyִ��5�cu)��-�p"P��c��5|i�e��2{q摥���a錦Hd�M���~�����ix�)�C��۲i����޲=Uj/h�)%�q�_����pa1�~p��C+�E)�Q-����Nt��8|d|��	\���"+ɩ9���I`s��11��u\�Gt+f�eDJR�� �*j5Ƚo��o�z%P�[��Ͷ�7��h����S��������R�Ӯ���vу%�9���L���w��D=�z�0T�����CF��l3
Rۢ`T���xĶ¶(�⌾������@�G�hn?���#�O�8�5,�K(�J;��V���T�[eL�#摝ZAC���ޢ����y��UI��k�d3?���4M���M �Z���eʗ��Lp�s`�\����D�H�ql��B�_ͩ��
��.\Is��|��K@�K&A��. /��b ]��xG0��&�_�,K4��ɾD⽋a�/6hj�<�B٘���9��rm�L�O����x����D�)�Q<)>���Q��)�q\)�����A�X�sжF���w�1�(�?�����cx�I4�1t4�B��SԠ@~p���T��ޅq��~��є��©I(1�x�pq}���0�!&�$�cH���zj[a��PL����?��9
�4v�ђ�����ߨ1�Ņz���
���e�G�N.[ۅF%��\�5�7�NmX�S=�����N���*���4���Dz�`00FU�E��~%�r?"���fq@�Ϩ2(Ȅ�W,Z	�M���)��&;���!h�R��e�k�G�#s��$��ns �NqIa���.k�֑*�l����W�\K3�7`�@�m�w�5�L~XB��aP4����y��{��Z�.Q���[Ed�iCӀ
�+�n�~��"Զ���2v��P��bʪ��y� ?��K�Uި��%��.�i���h�8d,�,�[�*��<�:��g�ܖ�i�1�#�	�r�7b�'N�Q��{MXZj�nOr�Љ7]�`>�&���$-# ��ElH3�.-JiR����O�V��$�|���[E�r�h":(7�x/��|^��c��й��b�d�k����� �K����>�L�uP��W�	K-�עr��k=z�unw:2g�;y��X�U'�=��#ߖ[H��^� l�y�vNK1n� W��O�!��5<k&P������I)\�Yͩ����L���&���B�8��;���"�C�U����м��E#ͯ\�oO5�����Z��|urg����,E@SnPq��M���CB\���q�X�V�s;@/聯K�^��69���<�fE�7Y�I�	�z�4�c�}$	ܙ�~u����G���G��e������@@��52��Y��7���*�)7�Y�mÝe���h�4°B����0�v/��V��T梜�=!A�(l8�<��̡���둈��BN�/�LD�S�%��] �p��U$PXJ��`�Ds�	=^J�<к(Jk(f�l��؉�rksln�a�k�q<�Ub3�������I�9[�o��8�����U�MbO(��&��\�b�m�����ukWg��O�~i�n�����f������ヺ^�?���:��.�z��?+�R+��'��җ*���S4�>'(��0�7��[�'����(����`�X�Q)��rX��4�7' \^�9������Xd,~i�2��B~���B�ASz )zZ��0�����2ּOn��xS��Grא��6����C�W����ht�V$�mI�ܹ���U/y��>{A�i�o],�J0n̴���vd�vpE�ʞ��ઝ�[���GԈ�m��Y��U�W��5�]!Ű�"����G8D��1�
��U��!��[<R��%-��u�KQiF��Ŗ2�ΨB��;N��� 1�c���x3��S��v����=芟'w�.�ʣ�i�]�%�G�R6���m.~�O��z93�~��W7И��Jo�cZ#v��W)�^k@Bm�L#�̈��.gS���<�@o��B�=�)�3�����/`{�0tK��7b��G*;�$S�'R�����Z�������
���H
@~�/���/�s�[ �H��_	2RN�`�\aB,s�3��y�<��]&�WȒ���ekc���,ߌ�&���5>������x�����zzq��ܻ�F���M}IGnɬ\k�A���v�Sڿ�Z�)��c���̆"���TI>xmu�Z��X"�0eh�NT�*YJO�{�Cn���B�L3[C)0��E#���<l^����M��q�1U� ��������/����]ٸ4 {�YA�n�>c���q	��nag �N+t�x��#o�a��U��u?�����ER�d��9�Ϟte��� uu]�L��,K��N�M�Kβ�^:�鼂u�o�פM��L=�/�� �M/�*3j��F���/ X
I�ɁI�Hj	�2�1����{���J����"�_�$�z��dH�ئ��$5G%�tC�Qʴgh�){'�����H���%�$�I���O����yl m��b�D����qV���Sl�Ƈ��VMz�D~�g{�	j\B��-�P]ǔN`�&#�9J�7c�7��3Xc����-ڊ������`�V [�H���[� ��*��������68{�R�v�P^Q5?���<����"��	8E�>�+�	Q�}𻀆6F������#~@$*�:�Ue]���М�-�T~#��@�M�@��6�]�M<����*��>��8Ŗ�������f&r��~=����$�˪{k�Z���.�����=��Y��\�MhI�hT�S����.�'���>��e��)�Q 0�E�����\g/�:Ə���2wX�Z�6�K���x,��0�X]E�(8������+@�\܌�R�ui����G���n.�iQ�߽��B�����I8���ܩ�v=�`���+,�k!E�*�<�?�����|��c<�}�����塑�V��L1����&p���j�_;���'jۄ%>���� �Gr��(RG�İ��{!�1�U7�ZM �z\�+����ߣ0:�`oS"-\ۤ�7z�YXwì�	!�P(��.�?;�y8��YL�o*X9�˵� *��`4�Q����X�6��b�M��)鐩;�	�ߑ���y��mP��&����%�E��D����ƴ�5T��Q��4CQ�'�-�sI�a�1��_���9~a�@�tEI���y�����M�@�!G�GL[�W������[��8X.�Q��.�������q)�҇�2��z�����9֣���n�p(����s>U�>�lA^
J����Κ �	R�2�3~7#����mIԄ��.L^i[����r�-Ռ:�Q�BN�˼Z0C�9@D Dxqܣxy�Oi�ώ�8���U`�o	5��V?V�Fx���H����S�j�f;x���#^�S���2�,�-O�#G�k#�]�Qk]�eKe_CP�qh`����B�s�Q�]"�|�����������G��زl���C*l.�������,�b#����=A	I�����x!l��"� t�����n)ޢh�PJ�Α�fզ! d���ݟf��]p��=��~M���F�{Zc(���h@�u��QC���2�C�f+]�� #(i|z�I��X �a��8!4dA�Ќi�p��M�����]��n��N �)�2����l��!�Z 5������U��Qr����XN�cְnhY�6����������f��U���ȅv_�aDs[xŉ˰=fM�w��ʷ��Q1����B��Ng�5������Q8��8��ޝ�U�Rp�o��
��~��gk�kQC}h�V	��#��Ѯt�์�D_�̛��}�ku�x&��1w�.������(<��u�Xo0QqI���h]������M�A��new�K܌?m`����� �~�R>h'q�SY	�קI��;bS����V�eb��ٜR	�s�!Ɇ�|��
�T\�/Q�-@ #N����
2�j%l����뒷Vk��_��tηD�+�迻�"6���p\���*5_CCW���`�/��h��΍��s:wG�nߞ���M�����|K�� �.@��������Ҽɸ*�����j�}��ͤ���J����(�T�k����5��-�.��:�.6og@�#��8Z�������]V��!�2���3H��4�M�^=o+)� �xL9~�R������W�%�}��8WՈZG�.��9��U���t9 ��;��8�[�Yܯ�L�=/eJ�[�J�KI��8�-"2���V�v����U(��- ��Bvc���%�\����)ҥn��Ⱥ����#^����������W=�}���˗=l��e1|,��'<�Y�I]�;�d~C�ҥ+yzۋ�Uy�R7����ȃ[.�������2%nV�j�:BU��=s\6�^i���vxϝ��:��==?Fd,�D����;ӝN�s�.|v�*Lnc������	o��:-��n:�ᑵrf���
]�ӱ6K�8iъZ���!b�!xg�@\�0jS�0��FX&P�Q�{`��Rh�T���[2^
Al�$4�V���Cs�^)񲒍����AENW^�{��)5/��gK�4���ݷ�eGN�a.3g�HU�/	S8X����_�2gqvT�� s=\���QG��]��@�Nr@���qYNZ�[�1u�l�p�P����,��dEp�mc������Øn(��%����W��R��BjZ��j���Bk։��DA�풼a�(�wC���HE��ɪ��U�)$�ڀnk���6)7��h!V#>�@Z����Ѭ�w���ǡ�1�@���������0������\e�#e<��&a(��l^�0�u�]t�F�c-8M���b���V�u�+j�)?�!�{�,aRn����.�1��zR]prf~A��@����x��������q�FE�����J��|�ˍ�q�n�K�΂�⢷�3���gF.KrË�@�ꗍ�k�U�1�p�'�.h����.Mׁ�Ňh1"�r���ʬ�#E�5\��"0�mS%��z9J{*Q1�H�o4U�l�Wv��ƚ�����B�"eU���۟��o��ڔ�'$a~�\�Ȯ�����b�� �'t>��$u��N1]ӭ�����A��"ry��"ϝ��e�лe��|�O�ů=(sm�e?��^ #!1���"Pֵ��Y�'�n̡�XZ�5`���$�5j$��1��*��|X��v�ޟ��D��TM��o:j@rhw�T��'ӳ���EP�K#f2.���.ҵ����IO>���OE��\�è^l�"�u5�LRT���/�h�SJϼ+i�e��'QTn���.'����n���O�����Pvҋ��]�&ie���ieIoMh)�� Y
���-��$ɦ�Th"�N\�D��h�6�K�`�n�b�*lT��2���I�\�@U����2d�t[��N���F�9#�*��`�z�*81��	#e��'�O��T�x�Ju2-8�7ܔS�!��͋���ِN7���cV�.~C(��7_�a���4tYҰ�!���P��<�G�T�|�5��Uy����x�h8�#�ƍ�J�!��w}̭u�� TQ�e���?�,F)^�'@�JZ���-���7%�}$����Oq?#���@Nlq�2Ȃ���[�7�N>mg�)׭"�g"��.�m-ਧXB���g���~�w��j\��2Q�㫎��r`�O�1�Ɗd�����ܕ��M����*�5�^�K"5��/�3�Vm��t bh��
{rp��>rzmM�?:5���R\��`��U4F��c�c�;&�v|K5�"Vz<��#����;���[{5��b^����z���x�.F�L�q�t���e/#5�Kc�ۑR!;���#Z�෠�X��f�q��8�h�Z�~/��ٳp��k�n۫HV��#�L��`����\����7����ǦEob�ce���݆��v�Q,`�4��vM�5Q!�]��J=����d]�]���C���"5�3��u��	X@4l,�!�"_���P��]�sQ(���j�_�X/�8K��Ԗ�!���@}�8��K��e->�8��.��<e � �m�}�'x&��f�I-�U�\M�_m�)t��-xht~��t+4���'݃:�>���N�0���� ��.���J� ���k5[P9ayWk�W/��l-�xB�3��}�Jm.Ԇ�TE`���&iB�Ϛ+-Rpԛ�)"�Mq��� ��.���؄���ym�R��Y�:�_̼6��څ+ܰ��J�!�5��O,�D(w�h������cZ�����g�o���a��nI|�?���rԜ�;+_mm�Cg�X�-����P>Uw�(v����͠g�t��W�ۀ������G�~Q�t���X7;�ِ-�A,Ide	�����ھJ��%��w9���D�u`�O��S���8ކH�~U"��z��i�=/�)��Ö6���ʞ|����G6^�]�|N�{5Kٝ�c<�	�;e?2��g�m���1��_��`@j�Յ:Q��7��Dl�����	�\:s��ބpGڲ_���9t''��o�bڌ�`X)M�=�3i�����@����]5�����=!�/E_Ѩ��}�U�Q/��/ԟV٠��'\w��x������9��+p�Ւ%���`y���c��l���qaJ{d�'ag��7�Q�x���ᶐ�(�徏��L�/���Pא�7�*�O
9�-T6,"�7��<P^00�dv,��^�}YJ�Q�ݒ[�~ɮA���&�e�E �g�&�-@%��P�/༃��)^�����g%��I&�ҨO
?���b�>����?�D&��U��YS@By�J���e�{n@�=�=ЌPaj�{0�tۤ��j$�j��0�B6)N�aC�ǟa�<�p���xa�̻���]����p���?a��/wk=pfٞ�
��T��=8�m}��vy����P�So��iU~�2͒G/�2����zz�\�ic5Q��'�B�a�{�;k�	��q��9�9G���3�LT"7��k��mx0��:�S������Uk8^���������c+�D���T�k��Q�PP�)�=+�L��4��b�)
�ˀ7��M9��~�M�`�p[�I��)฿[=Z
��ȥ%xG������V~�n��S���P��ys�b��'�H%�LHThe��]�!RG�Ĭ�m��uu��4Y St���c�vJ���2�5��$ǐ=s��ꮃ~�څ��P���2�O�%/,ɦǘW�Z*�/$�7�Z�ףz���֠���[]��y�eR	\�`�yI� �hx9^�҃�3򓰍TD"�Eucz)����r�Ú� *�a{~��S�$p�^��b/+$ٽ㎫�ȳ���a!�f����$��"\�e^��qz|	ʦ$�`I���kV�c���f���pE��-B�₼��.���H�*�%%�2��C��+"B���� ���9�,��e�V�5�B���y�g_3C�TS)��۪��l�ے~o���F�*?�><akz�-f��#����Վ;�;�-RN۵�����o�}RVe.תߔ}VΑ��	fu��|�( M��Q�|UԞ+����������w@Qr&�}��o[z��	�J��=�&��^HIӯ)5 &�>2�k� ��>I�D*[u�"�nT�ܬ�Щ|�)���:�P&����4NV�UX�p����
�v%��T�LN���M��ꋕ�4�1Sˌ�.:
ԟ�#ƾ�Υ+������l5�����(fRk΀�N�����7?>zCU=��3*G�N _��O:7�2���kI`�;�q�C�f�>3&�D���*��3�V�%��=�P��;_��1H��D�o-͢f�l\���	�Ơ�.GMm+�0Ly"2|�3c�����rh�i2y��}#�ơF�pL�*�.�E��?'ůXa7niw3:s긃�R�I�y��;�$=�l9�{��X{�@+��s=�y��σ΄���3�Tr��	�}�r������|x���$�K�m����mU�@n�G�4K�ǎo9BYB�7U1P����b�mtj�>X���JO�[����WE͉��-�ْ��ݹz⢨<m�P��+���n�/H�5�T�>�A��Q��ʛ-��.3nu���-I���>CΣ�Bǳ�f8��n{C�QY����c��t�A8��Ѽ��oD�iڣ�Š��[.^�;��w�J��֘��3{�}��䛌��Ҙ�؜�,."��5�Hm�:��&_���W���S�wƩ��{a4y�v����)�"K%T_۔��N�Al~����lGNC��[j�9���*|EaZ��@������id�k���~��P1v ��`c+����(���f��ax�K<5Q�Ev����ַ�GK��H�z8�b�o���sqw�
��mw��t�������3�X4pD���ϗ"t}���4�3�.ϣ̊�Ի���C/9V'���%�����(w��D8���+:IQ�GG؏_I;������v� ݏ�&5my��䂭W��;/w*+�!��:��r}}6tn�M�M%�m㻊�ۋ�4	�׺���Ⱥ� h����?��;�m�#�ݿ&�̥:^c��I>�N�0�)
��_~JNW~��k 	+�����x6��KO��6K�3�M�aM��'�&�H����dYw�f�Ƭ#b��jMo�@S38b��#��9�ȱ�G"���!0
���A9$f�`HgJ�����f��g]���fB��F�?ҫ�׬-<��z~�C�!���m�{ �m�~07l�����y����9������۶����6M��4�>��r��l�!��5�)ر�<�m����_���J�^r�B�<��|�N��2Z�H�Q���!�XЄ���y"��d �?��3����W�!��̇�RGfH��M61>	_���>�f����h��x:i�0�@@-M����[�n���㰽\���v�<�s]9����,��yH�L�@�����Ġ��:�
����Oa��R�)�������ȼ��wa����k����?�U�.���ٮAxiQ�^|iI����J�m��j�����*ȟ����~��{TI���%W������˞�7��0���)/������G`��AI�f[)Ą���I�K�W�]+SxM#1Z��X"�Z4�c��M6	��t�K�	<���B2�JӲ�����y\r�����>�v�q�cD�e�+68�$ю�F�w�Skjc�	�@�ē�"�:�'�9<|\��+��E�Ry>�x5��$�Q�����*}J�sR9w���<���c���}�
�E�����wn� �|R:.&�{�p�|>����Ô{`l���(�H����ER�D�J��@����g/�w��%�R}��B�H��z��M�$�2�e�ҝ�i�1���1�^���=y'���0F�*�o�~�u)�y]í�pw�C��6�pO�<<��(\�4�w��U1-HâGQq���s ;o��ŒIu���+�����5>	!�����'n��{>Ð��,���KZ��N� �	��W�J	�uViz[i���f��t�r6&ė u]��A�hO�N$Z����+�����s	գ���f���� IS^�Ƈ�p��j<3{��vH"�wC��\)�9���h���Y �W0y*ͭ�@(���J�O��s��^��?MGLH�
 W�S��K���E�E���O-�LB-9;oz��q�t��E���n�(���;��c[������/�u%�g�W���jW��k���Rj@J��˳m�Bp���gCqC�Wz Y�����q4�1��@��������.��Pu�v�̡K�!
G�O-�W�/l����ך�u��T�,�$\dQ,��v���P�_8��u����(xp�c��E~PP�G�R�큵nt����G��B�&�t`��Z�"�c��j*qn~�����I�{	��g��iӬ���dT��ǳC��NByf��5��} �e�G��"���):��U{��؁��k�O��K�{4N�[J0<�ͦ����(Cd��(��\�����	V�ۛJ�2F�^Gg�42��	/�6�JX]?�sC8e�1���=&���sh�s�)�1M�<�=y#�ު�T���}N��o���A�ۣc��Q��m4&�lX)@q3��0M��s`qz��D4��_����y�T��k�@���f
�]���8&�����IY�<�K�0���4�l^���[�^�>%�9!_�F!L6��dٲ� 	�=��Ù��:A+ayi�B*�L��p�����~9I��-�[��!P�+Q%�[��F~٧�� ���I���Q!xe{�ͦ�J����*���|(cm�Ȑ����x��U�9�����5�Ok�dU����5ĺ��;~ ɘ�QvI�L?�=�7���c�����P�WS2��>%�$^�Uu�%���#e�ܿ��d��"�p�&�QGXu��$Z�_��j�i9��-a;�[T��v��˗pz��:]�TLB��<a�5�#�w�S�2
� g-E���!]�ƅ�}K�4�Z'xm[a.k���W3#DQ�Gg7V�`�}Y�ܯ7_�$籜@�#�$z^����2��mP�+�ws鯺��[�"�󳩗���P"M���?�5XciʦU;_��8���y�������a���%Mu�o��C.�jO$�d��:X����9Ƶl������p�P!F �Z9�xW�K��:��3�?�a�  �xj�VsCJڛ��|��r�^�1����z�Ll��R���<c�/�8x�'�H�u��II��<�%��D�ˆ�cQaS�9ecP�yT����8lu1ٻ���U�GOgb���J�MK@����l�׉�c<�1RjF�]*Ba?�v��4QR��%7��o=Q��N�#A�E�*`��^U���#�:.��϶
6{���� ��=(���§8/»%�Վ�l弐_��g���,AcEKX�?;u��X�õ��5AX�c |�~�&���5�Ef��vN"�+�ۓ��j���+�CJ4���gJ~�]5:7R����w�f�ӱu�8�%�[\O��d^��-Wbh(p�	;�����`	�1N����s��
��tӁ�������8�:5<�m���ԆWm�Χ�U�0����m��z#�|��:(��&�Tj�P�̼��7d��l���~2b5?\ W�jw�����L�%��pm<��*1�L� (��L�)�d�D����&}ʋ�nӫ������i���w�ihg#���̬���C$M�~4�d?f�]m૸��y�z[�������9Mn�:���^:w���­X�m�	;8kr�﷯�7�;v	f@,񻞆TN��Ĝ���y݃jt���H���m��]�)��r���F>�� �D�E�o8U�؂S��}�Y5۬=sp��G�Z��5���WEn�_5�F2�^�V����%�H��x�����O�����>�y����#���Ɵb1ݐ�����J4����=�K͞��x[g��W�р���$1��q�ܭ:FC�7������E�i	�.�#]��z�r�.4�' 1]��iLJ_�6D���0��惔���1�9�J,q�$m��ECB2�P�+�����lTmf �=��ޯ��=��>�cu�����1 /\o����G{b�ʳ�%�"����{�^H9��6�����XT5mָ�������ә�W�����z�,�5J�
��&R��/�����[�&�C�����va�{������I�[�Wį�G{y�װ]_��r��2�T�'������߲zw�zF홬]+�Saw�U�bQ"7n�[�ab�R3݅;@�H���^5�E5��4�\14.����kU�����o䓺NIyʇ<�f���4��I}��h1B�>�5��T���dƮ��ݙ_+Df{ӹ�߇�}>6[��/k�J�8��?�<�82���$�ޘ8Cps��e�64괒�[H����3b@��n\^NU�+�O�f��U�S�.BB������iؑ�Z�� 6��q��ŅϨa�f�s�bO�=��AB����4���"G�})4���iasW�/2CH�1�# ό ᆦ�K���R:@ټ�Z�(�U�t\�h�fƯv�0$��/��T묬�D�B:sm�x��fm��F�=�(G���j�����s�g�q@�C`�%|}e�ơ7�,�\��QzV���d����?���k���|�b�	0�D�>�n����$�\�,��%�2F��,�n���p.�Y�ua��"&u��������;Su�� `&��68�pj	��A>7���l���� ���R4]T��u�w0c���K�M�W��IZ=�4!� �fh��Cb���@�q�z�^#�d(_�v�#zu����m�pG�n���0���ҌUL���/0�����vc��m�3��3gH�(���jpwC|^��ԯG�����܅�R�nG�$?" �ryxb�����v�2U�	�� �������p��O��®�Lt�*�;P�N���1J=��dH�ͦ������H������Wp���D�L�:��I�UG��k��׋vrۏt��0�˗�(�f>x���a�4�k�݄�8��t����;��رb��+ !�ZDaӇt���Ή�F�/�*EX8�7��>��e΀2�М������ټ�^�/�S|>�q�0�JA'"lcǫ�������H��,�����ٴ�Dɰ�����[���Eu�����	 -tOkC�
�����mۜ�rgc� �^��^�9��qd�Pn�~s&�G{<IVbE=D�Ǫ�2�u�� ^[I���~"�QW���!����᤬QQ SB1�q<��U����|$�"F�̰W4� :�h�������1���9��Z]�`�� �uډO���(����o�T{�f�	Z��Ε�}!gc�I���y%�j�w\_[�*yCC���R�8���@��&4�RdqJ�tvA�8��q�ͤ� E�!?��f�#����\��e��+��fn寎`�P&t�c��wa���͟���IWd��y�ð{a��>H�̦%�R�64�A}�1���o��f	�<VA�;��W�j�C�����g�_mX�E��U����_Br���(��k�E�Q�^x���N�o�é`���~:��z�!_���|�=��p
@.�y���-T�V0�VnZ���I�L8D�4Ŕ�N�n�3�&���̤o��klY��r~yͪ����YT)�6�`=���D��!XK��,����/~�n6����z%�wē�*�������
�6j1��o��A�ȼi-�@�3������|���WJW+�y�����N�^�����Sf�pu�0� ��!j)�V=Q��:y�w䅤���m�G���np�bs�A�����i���{�9JD�?�g;��AF�Cm�E��o?��?uu��S��A]�h<1���!�� �C_�����J��7W(�I��nf�%���F<�2�X kp�T�w�YOCm�N��5�[��IJ�ܶ<��z/��[�~-He�&)�+��L���G֬��,����X�ReYө��<I��V�v�g�cW��~ٙ��$��S�#A`�R�	D�U(��&ܰ��V�B��q�v}���(Z�(��Zw5�B�7~��2���J�� T'��(��f/���_�%t5��4#7b |���_9����1k5�����HjI�a���#)�N������$�1�b�Q�a���\�e'ˈS�Mvd�כ𘲢�s�a�l���)?���{��̈́�ͥoz�	2
�C_��������>O$yKXw��鸞V&�8K W(�4�p���D��q�gMP��{�k�����ac�.L�N(�׼�1G<~)D%:�p1Ս3I +m��E \����	�Z!i�O����'��UGN���t�,�=K�/D�A�������<�I� 8}R)��~�����.\��T��^�-0=Iڻ}*��E9��~n���ٌ�+K���� CEb�&�	XT���"l!��ʅ���c��t઩Tj��
�͞���� �Q���B���Z �C�5l���/�<�L�2���kŻu�4�Tw�}b��lUǆ|�z�"q&�B�5~������^��AAQ����+�\@wA�L<d�xa H���_`�w^\�����<��@>5�p��� l����-:�����S����K�����ۑD=�ϼɮR��m�7��ѓ@�3��K駆���<n`2�()�neuQM�Kdy��T�l9B�5��!>��o�8<lS�������I��ĉ��� �@3[�(Fp���u۪=��*	~IO�H�k>��RT+��طǽ���}$vDnm�'��i�V��,bY�g� ��WK�X�a5��:���	�2��<A -��U�I�1)xҘ0M���1DF8Ƚ�+����+79D����Oݔ�3�[D��h:	E��dk@�M������5T���|��jC�	��3��E>Uə�<�g}����+:�8����8,B9BI�g�'ˡ��S���KC*�]�����d6h3e{[�$�B9�f1�iU���9���\Ò%Qv���|	�����k�X�O��0Q��e�ɖ�%T���t�T$��涜�	a!�${g>�>I8w��^�O�y�BEM5V�.r}"��� �i�ѕ�UE�jnur�{�	+!�W�zg~H�:'�-~���� �~]��I���Bx��ݩV���k���uY;�@�8�%��	bFD�����\��3>ݧ����r�4�U��r�.m����]_�Y�&J���|�{">���G��CA���Ӿ��]�W�A,:��D;g���۩�i��Hf�5,��z(�Pu��!i!$�/�.䆊�����7:FT��3��=$����iB��nY���	�զ/e-�ґ�5�)�u����i�e.k뺂�_�O��1��p�K�����%�x�G/�������wG'���^���WOK�If@��Q���!M�meC�6�X!L�mz�<�
	�Y�G������* L�Ws��P<�24g篇
 �<.�qs��a�Cܟ���h�{���݉T�҈�-�w~�����j�Fxk��b�|��;;M�> ��Z=vN�}ZwKe��z�tz�<��_� ���~�$�|C;��#`�U��
M����e�Y�:�b�.i���������[�v�v榤J�P����\��b��b/Crn�Z_�w�9�v���)�Bl�P0���(/!���RJI�d��YEʵ,P�#cO���V�M�A5aQN����y��I"���Ec~-��~���� ��'P�q2 u홳U"P^����ց�I]ܜ�+���p �H��N�/:y�Z"2G� � kr�a� ��WjHf��e���O�p�T7��:@*�\���*�%M�k�k��j�o:�~#��B���RF-^@�@�/F�AK*G!����<Cx�HȚϢ� ��Ы�Y��Y�8��K)�/�)J��������Z�>�7to8+���ee�??Ք9pI�'1w;��x��FSǔK�iܳ��dut���R3Xi�G�ޣ����L@�i��(x#�G��W�^E%�N󩠤]U�T��mi�+�v��U��M�]۱ɜ�Vp ca�'�0����~�J^Pأ�lp t�|��H��lm��@�����B�@$��|�`+%�V�Fv8��	�
���\m�W��(�.��˰b[@�C�Z�Y>9?�ү��z�Gb"\/����e7C�6쑁�e��K)x���0L@0L��'�.��l�g�oy,��}�s` �{��9����0켯�^� ��!�-}�:N��y��n�(wn�[F4d���8�$�q��j�	,��	��x��88k )����HO!m�]�rS	�27���G��p2#��:`�X}����J�2�Ϧ��=���p�j�{"�E�=��!�Kj�v8�y(-�S�0|J��2k��*(���@�m�ȸ��m�w�B�7�Ʀd��$u jb��JnQ�*�n�Y]��9�;"F��wʹt�ݘ��$�{��Y���}�6� od��Sm�=x.�N���~�Z܄�dN�����j�_)�A�C��]�Y�%?�HV�8�Mv�����N���-�5t�:-* ��$���r�� ��e��qrC��|C$�3�� ��M�D��YE'�4�î�y��'Јǣ=�a֒TSp��ӜشHO`� ־��h���	��+�P�W�I�|�O+�>c��Wf+�~}JA�Q��J��6��^_��m	7�_�%VVN�50R��q�r�7r���y�;�:�عYKr�R��#��z|ѫ���Y��]r2]\��'��E��i���Z���Y��r�a�8�)�+@��}��
��Ϛ���p�@*��e���6��̹��0m��x9������p�o����	ʹ�Z��b��O�q�~N��W��L��z����1h��
��GT�9�ݍu,`�ߴ��Y�b�4b�W����ӳ?��]J{��^J���?\W"��a�
~����(3mLM����C�ݕiV����9�_ӓ��fm��,B�ov�L�+[}֫�b*�����5�T27��p� ���uF�~���;�B�*/�֬���4� �Ę���':m�B�����Z	)�|��%۩�M0Y��*A�\��7�z�I�!�\V���Z!{Se���a����;J��5M��|�S�)@꫻�/�dmS�!*쀞��a`6�(�O|�l����':�����h�jqd	�J���������1�{AGjw�C�Mg�P�3�\��A�/���������;��-k��--�9�.ҫ�ߧxJcp�����n=ˣ�m�k=��ִv��d�tՔ��6�hB%��9�E@ڪ���vVEK|i�f���л��7���v�ہ��=�d���e���X��sx����IԽ�Y"�zV��g������\�^&<.��f���2��������r�"�B�z�~#���P����ǔ�G��޾�s瑍�P�S�곌ha�Վg���wV�H���C�f�H`��"o"�|�_��;	������Ӵ���6��P���JqŴ:Q�  yN�R+3�4�G^i⼀6C�A�mE.V�;ƹ��A��uBRx�o/-���*�}��ԩ(����-��&�U�d�O_h��\��5ezk]А�@�+�9EY&\O���;��Xj�_Tw$��u��!�&8aS��`,w|)�R�ǿ�- �~f2����A��U�>qppP�(m;jk��V���u���b
�^� � �U�8���44ܝo���T�z�\0���ɟؠؓr�ɿ��W�h��x����y��!�vny���;�kK!�s_m�Љ������Z��t�
��[���pq���>�V�����+{H[�M���&���V:�m0U6�Va#5i�k��7z�z��my�q�A̹��J���Յ�n���+7���9J&��_���}hAƯ@�r29��t�.;�"�.��.H=uá�$�$��p��^����J�F��Ρ��x� ��P��*ya������n�y����p��79��GC��5F-2����uSc��`[RH�g�ߺ(�JS��"�"�|סd��,�W�:	/ �#4�m��<�����Z�lX�a���͚�>���'���jz�_�z7"՟�0��P5�v�+����*[��ü�a��r&W��r,��CBE���vD����[�uUN��R[k�k8$�����FB}�ymZ���P���ct�ʫ�B� �O�I�P C��79��!\��!�.0k�
I���t�*��A��$x��[LԬW�5/a'���p�V����u"X��2����]S}��[���b\	�xVnI���
"NdE�ivh]�����9!t�8싋8/eg���Ƭ
�Uw�5	����1�Br���<�~�n��2ۘ$5�֕ܫ���`'���#�]D�5�؍�(�m,26��11��`@�m�Q�vf�� Zܐ�2U��W9��}L�:�	��M@Z(�W΋�0cѲA���j1��0fF��]���x�A��j�dg����c[��V³��Z�^�Nݍpd�����F�h�q��#l�¿��!/�>�NcG̞1o����ڋ�,0&���L*���{Z� ��RE�����:�U��H�4JhL�X�!`�p����ފ�la}Al�^|�9������n�d��0m�? ��\����Kj�lm �Ex��E!�w���L�K�'�Is�0˾lS0���b��ߙ-Y���L�jSR�Qf���	�3�m���˨���_����7p���Y�~p�z�"�Xr=u���^�S���!i�Ig���v_�/Uj@�M�q�HACS��}. SH�Q�E�~-�x�o�H���f='p͔�v錂tc���f�x��?۽M����Ѵ�{U�L�ͧ�(B�"���bJb���`Er\�FܯB���zn����*�}�=	1��Gθ����1O��r��Y�R(�3/�S��~o	��-b�k�9?Ը"v�6n�X�!XWՒ�ٚ0��3�jW��V���-áD�}���L��n@4(�Ɓ`�jh��?�)rgPJ��|�##%��Y' og�`�@۪�o��qe1}]��RbOޭ�3�ZNN
�N?�/�_=�ҥ
�@�:�\`����-,�{ �Q��}W���	jC�C������Ҝ��Gkc����Q�L�9<��J�-�):�K��ȫ܍|Y����9�+�U�+(7o��.�>B��H�;��غ�\7[�y��n�D��D �{�����^�An�QY�������j�z�[]�b����D�BT?��"L��&���Ec��ʝ�X�;�hpI�����Ug��C��ڭ<G�¬��s^�6�<�H�]��-��C�GK���A��G�j�)A�-)�IR 3ë�>u�,�{�ه�/Y_554c:p�`���'�j��uս�MK�|ɽ�������A����_��c�WM&�L,c>@�߁5s�2�=�ʧW�{��Is�%
a�*j�z�'"���! ��dt��

~ֻ5�B����R�_E��Z���~�#(⥂+#�o�*�^��z��w�D`��/
�h��Ka%�}&
�k9���|�
�<@b�3;�m��bk��G��zВ�
$�flN�MD�8"��)�VO�d�.��LOP���B��@���`���`�!��vn?w}f;cש	��ׁ'�H�<�fO���y���"_����zM�|I=v@����ǁ	�y�v�-�E7�����݉�{ƥb!%��P"&�	��t��+Rٗk�(��������V���#}���Z��:�T�b
�_�^U���uH�8׸�6����y��C/(���3s���BY=��+mGy��OX:>g ���n�����w#�R�a��^Wӓ�&�S�H ���L6�Z���	����%Y��F�g�y/� թ�^,����c%����-\w�	�B�RP�6���)���s�	r��ߐ��QV�+�fưN����savL��AQ��b��V�6V$����'�!���m��G6Ye�~J���&��&x����8F�-�R_l��1x+������y#�n�w���G�ty���݉�����%�K���~PND��D%@D���e�G����jw�~�574,	�S��]���R�����z��(�y+���
��Ҳ�Uh�8ot�9}��b%O��Zcٚב�曡)�f.��3(�xL;*�����I��HH5�G5�mHL���N0��;��}�0j+f������5���ec5�]��;��	7.)e�&�˸a��/� -
n�l�����b�u#t�Z�*��2b�{V����X5�5֏�W_�')�U7(���Ƀ�;��5i�6�Θ[��%�E�]r�#Qu����,�1-����ٕ�@W����sQ�K��gk�I��a_��L�U-��8�D7$�L7�������̵v�j��&�P-�c�ei�i�5G�-�˜�/����u�����3u�5Օ|�� ��I��A�_�Ln�t8��f	�f؝ D��*��A�lx�K[x��!
������j�y���$p���+�=�����.]Z�����5O�Fi%��o�2$iX�� u�������f!�����A70�@��VW� ��&�M����6'������;�J������]U��pZ*�,�����#72pM`!J:8�6t
���/��������Q����0��Y+qY��E�+��D�	���}.�V=v��O��Y��D�-9������\��>>N���P$�!���j\C�_�������*�o��Q#>�>���c!�	�3��9P�?������ޟ5�GZ(���S"y���q��0ʎ�Y4��/	��ZQ�r�S��w����: 3�M)�nd�Xp'�f�G�FC��hp��`�V�:�QX㥭�e��zFQ�E9�K��ų{w���ƣ���c�3���[3���2�@��}��d�:�8h�02o�T|�R;��)i~Z$K�#3��v/��"'�$�w��fQ2�i��T�津6ƞZj�x��[�{��^O5sɕ�� �1+���৵7Q#(�i�j<���?>�Q	0����|}�W$cC^ɀ��rm�Cu`���9�űv'�L�M�q8�p��l\e�s�1>2؆��)�4<�j�ry8w��+�~�l�h"�0�$9{H�lh� �eu�w�GP'`���Ƅ�צ[u�y��J�@G����-Ҡ�K�S믡�%QknՐ+27Ы��W�r�%c��?�r:��B~m��N[��)�%.Ci�y��9�xd��t
agH��3�,�$�摳�z���X_,��#{lc����O�����ԫ_����Adk��i"N�� �����h�EE�ڨ�I(f��d�5�NÎ ����Yd��L͡X���r�AZ�x�}i�#�#�����BE%��ì0����}�Pk���jȣYƷ����WE��yL��ɀO�'��8o�^���m���]�Ç��ט�_��Ի�1�~����ы��C��^�#�y}B`Q,��.Jި�J����U�Q�)�����#��|���NdM�R��UrI��0t�L�z	#.�a�K�C�W7���{��P�����	�%��xr�2y��������燊�:B���\W�5��њ$�nB���U�g�>|��H�4�-�࿍�ӻW)�'C(���
5m��K�W�ܶO�A#��y���(��	ޒ�֚�@=�5j(���h����"t��["�7�c>���
��y*�ϛ�6�,���s�\@�#��0���k��mIQđ���x�Ou�n2�5��3a�3��}aa����W�Ͳ<L{j����]L&鮐�˛�03�_�"���Kk��0�v Dk��jۧ���e2�� ّቬI��8v�x,�S�?6�x��.\q~J�g�dt0�`��sڋ�]E�`����C�_x��v��Ju�9����-�q�[�곙0~m�E�hm��%n�!,L��J�粰�n&��)ڳM�d��n3��N AG#�_�l	�̀���.� ��N���D!�[��pt�k>��l��:j�Rcָt�N�.�|�3S��bi줂��g�.�1��#lt6[y���O���ngy�~��^��ŹSy����4�:����5O��Ib���%��>}1 �C��Mص[lcဎ��uJ��? Wf�L����AE�.�vf�1عM �~�u����͘�K������7ky����j'g싐��.�6�M*��8; ��ƴ�eF��1f&�f�6N�P�J����w�N�!��c2Jp�.��+m"����u2��è�OF.P���@������S���3*����q�瘄�a_�$|,�?�oz�� ܼ$E�e7s�*��iw'�����K�hv����}�1 2q��[7ɳ����@8O =~� �f��u��h��߿n@�~�S#!=�H�y�;���A���^&3҅		p��j�R�NQ٭.�Ήo���[�w^��m�8x�yE��wc�O������`��	 ��©��ύI5d�5��.ڍ���h�5�i�CDG�9]�g��/�'�	[��p犼DW$���E�mw���:LK��v��c	BYmY�vj�=�`�[|�����y�`�m��3G�?f����;'
Q���B�����Pǜl�9G��S��z\��$���Cr*jOuN9Ч�AL	{��=�9w�NX�+"kJh���"�sV9�:��`����>�b|mAA���M(.FAo��(Z���?��M�J�5��4��&Ly#�s���a�H���e&��%( �;�B�ԑS�d��m?\�� l�:��ś���Z�PY܌R 0�XF��U�^F�sɁ�t�`�|T��C�|dTI-��u�&iݶ�ՠ��< �'X��������&H�;jo}�ʨ^��+��F��j������	%U�����_Idɺ�(��_}��'V�G�Ց'�BO�%* ���Fc�wB��>��H��r��"Q��-�,H��/��������F� ��1o75�ͩ�,1fx�˿��I�X���6�uȒr�����Ub߽.&�/�H>�֢��}c��p��˘��
��WZ����7s����ac�Es��f�|6��e�F4ے�����ck�	��ₗ�g=Փ�/uDV��[�!"nB��Z��$�8�瘨�� q
����[���i��s]����r�`3�qƥs�T5��Q2��da����kf}%@��E��v4������_����H�[5U��ѓ���qo<|��'S,�1���,�7�IEz�l�|�"a��Ϝ�F.j��̊��i$]��U!�Ϗ�"�Zz,�4G��ω���[+�y����$����R��;��Mybj8S�8sF�7<��ǱL,/@C�r�>��Úv=�H�%~��i�0�R�;��l%>��M*H��L]k$�#�����m4ҹ�v_��%��vq��ڐlC
�X�&1�6�wk��N�6�,�L���
[v�#E^B+��I:�2p��Q�R~Q
�Y�K����d����y0����G�W�^���_�L�?���Y���u1+U���|���<��ď��3��f%Z*�O�Re��f�V���5�H�4�!V@���"
S�}V�D���q�|�9��*
T�%��d�Ǝ��,�����50���ޥ�Ң��[�Ip̟of�00��ꏊkϝ������M�ډH]�D�gH
#�.�3c�Ɇ��i�ש��\Pl���ۇ���q�HE�0������s���!�6+z�_��9�M0/ J���
n�	�c��ǒ�Ć,�t��qN�����s�����~��, y��l��i(��������3�m^�B2���1s�4ⒻO��no��u���P���iZ~^�c
�	��E���%!�F�u�8+S���(q�"Ui@�~Q[�T�H��&L��)7�N+����x���\4�#���nX#�&n��kJ� ˙D#��#Ut�N�.RB�4ȸEv�eh3{Oݟs�L[,�*L�L?���9�?�՟I`��O���]�C��\�&�k(_H�eDd��8[|��f;!G�W�`z�I�k;;��3o�8����S&��\��fZ2��߹[�|�����;�AL�@ZY�uj���\��^���x/���>B��[���]Ш���q�(U@��$n�I��W3�JTF�������
��T�0C���������]	/���a��b����7���^Sm[�ڤ�	�b�L�/O/LK�F�s*�ΐ��<�8�;EI���S�j�J:��D�8��m2v�4�W�����i'MQb���Iɕ�b0��Q&\��#�G�鼽AQ:�P�\O_��u\z��C��J/�u���^�7x ���ļF�>�(F�E4v�mB��>x�d�|=�*S�`g ��ѩ1���(݈��`k��Zy��J���!�7_{W)���i�a�js�;���;�����!���D�%�M����(*p�@�D<�Tj(5����e�Y:c�sY�p��"�,�x�s�~<�߶j��sb�X|ZG��D��d�y����?�5Xs}Y���3�lC�h�^��G�s�ÛӶ���$|��%�/��Lo����^4�݄�Dz�����o�v�42���b�$o-�G{{QqIl	v#�L�t|>h�����>f~����P+�_���rNr>f�ߣˀ!�{W��F�<3�q���
��B���J,��|bwyl|�ݼ��.K��"�&8��f�6T��f�3��L�J�P4[U�D.I ������->Z�k�b�a���J^p�#� ���1��0Q>���گkR�_K�f�6N
s �ޒ�&�t�o=o�+!���f0j�b�9��pWd�Z�"��+u�l=�}*}��:ҍ�L�3�
�8%}v��ءe;\]0%h�A�-�E�?즲�!��Ծ!����>M.�P����a����#���5�'P,�)�_8�cu�t�lb.��c��p�q۳-T��"�B��dΜ]�H��d��2m�J@s�}k���8��>�͛��qr
�0�u@y�Ź�*S�o����-Ύ���X㌛.���!�iԣ�GV�D-!��IWj;��a�Jn]Z{�Rs���F�@K�_YR0�z�8dQ� ���4/!x��+k��Tsh$�ǁH7[����AӪ��T�����A"@���d��g\,|4r��޼a��F���Q6V����҇�X��JxT�Wz�G�ۺ8����o�~�_ra�4������&��|JK��n~��DW�|k�#�+㋁��#����4`�>�WrSP+�.S
�)�&�0n�2���-��G�~1XGw ��"�I
�g��D���bڮt�u	{�#���'w�Ҧl���P�u���/șP�������Jߊf�R�Tz�*|{�<��,탑���G01r'�{]�y�}�$X��)6˱���?4~�L� �j53��Ξ�]wj$x�IG��.�11�M��~��W
bʷ^��R�VڨG�;LR 	p�C���[rZ�T��HQ�����#���|�1X�޺��H-�$;��b����Ы]���퐭"�e�a��2���=p���mz� ��N#���})�Y�p�]�������S��C���a��MK]ǚl��q���iЉ��~���^�.	���8�8'hx�)A�����^vt(r�J��t5��7���|@2E���!�����2�U7��q��#�׭M{��_P���6��D��|C����{��i:�.Fj�G�*Ж�PZzQu-��I��T�Z�l0�(��v乗q˦Po��:�mr�:Ƙ-�NM�� ?�i�j�]�x��⋘fyQ�d�Z��B1�!��y0����'\��
j�Z��Ow�%P L���`ڻ븬��"�P�38����GM�4��nҰ�3(`O�)��$
��,D�O��W�W����Ct�T ��T+}�0�
E�ۂ�@�/�ț�Bbk}Kg��5�l�J*m���n�В��(��M�r7)+LtL�I��sl�;mg�%�K�`���5��7�w�f��GL=������u��n�sµ�g�Y,isl�^ρΨ������|���Gl�z�;'^5�����5�ZL��J�wƚr��y�k��R��I�^4�UÆ���
��b\c�v���%� �F܅�^�dJ�}���"��w�wA��K�5b�o�^�fǳ!ؼ搥�F��+��M֢���킺�ĂZ�H1���~�eΐ�r���6���'Y1�����t�*.�#~h̜k,�n̝�$�E�U�v��=�d��I��|u�>�{Q�m_�[�tDwrl���$���=���&S��S��@a���,��.=z��+��S�xnTm����B����/���R��|�	S흧���2H[����U�9a_���d�`g��a:�A�X�B7Ӻ7�ww��e����$���G��m1=�o!qLJ���J��t���4^�U�p�=՟ ���l��[��1v9����xCgBP��`����p��!u�4KPYB��5ϲ��������m�v�����E������E3��~/��/���b��.�� ���4�|��&��y��ſ�*'�rds
j�V�銦�i�]*%?�y\1!�_����aj�U�b�����u���q�Ty��%�{���vQ��q� �ΐ6[@z���Q
8���Q/�Ԋ�ɍ#��Ii� �%4rx80��g�u��"x��eGt�f�ߔ���Gg����9�\�z������7�q�2%��0�w�Z���z6nIA�5��}ε�y�G+\�#��):���8��J U{�P�q�5ܖ��1�������-$؝��ITl�����@M�]���?#�!�Q����.a�F�(�?�B;����B�J�����p�Tr�D'	�(x�5fܛ�|b����A���J<HBL7�2����) #�y!��f<�����5��r�*������p�F��S_R�Z�I��������$� ؤ�U,I� ���V�����6̫
 j8���#�ad�w�i�y\����7�n*j��3�b�o�V`q9~X#�#,�hFh��4�ږ��mQ����7U�g��+����(HԘ<l[�0��L� ����)��T�j�	�|�S����.�k�ϑ�^���ũ��NdSY�V.�7W�sߡc���B@'`��	�Ĩ��I�;JyHF���lQ� �G��~߂��U��4�L�'3��@-nq�G��m�yT�e%��
��/p>lW�'7�f�3�)���=)�G�4Qu����Ѿ�HJ�j�0���/��)K���w���YP���*{������j'[�m���
:4L)K'�lX�� �(�#��^��\A�R����L>kV�~��绘��9��^��Z���}P	gW�	�&R�-i,��ĥ-�i/`���RM�l�
��&G@�bGAi$W���i^'�U;���	�55j��_~�\$��Ì��Tl6��d����j�ް�Q�� \��Jq�}�9���=��M���┩�+"ʶp�b���t�������ʼ��焪�5���fr��q�r����(5Y6��e��@�$0��=>gj^�4i]j�?�ҧU����y��Ζ�Ɓ�z�
|}q6�����X?
�ߐO������u�����"aw%���0�S���Q�oW�;��:1�
u_9�_S��^m��cK������1E�q�V�������$��&�29����TO�ܸ��{�t�b�-���$�}߿T�S���/s��5=@�ؘ hYcltm7��Y	�|SzB����J�}Z-�<�mT㒓����P)���
�t�D�e�"�z��w��<�\�L���9#�F*"���� �H�6�T���S?F��B��=2�C���x�|y��?�E�O�𩠐b�r��R��G&����Fx��.�R��P�����{\��e���̺e3sQ��ҝM8Ci�7ka�F%��$��ɥ�4��?!�����3���Ű�I�49���8X��c�~7s�R��)#�x�Z�+ B�[w����2I���U�� L(��S���-R��)�
S-bf^�٥?�#��m��5gJ�΍�`�%YV�i�|��'��壓V$��$5`�c�N;�n�����1�͚F�3q]�?�>���JrzT��D����,�4�B���A��I��[����G�5"���k94�ss��CVӳ�^dB��q�v�0-���*T�V���(C髎��g�I����|[��@���ũ
&4����2�Q��������7{%D�Qo�a$VT���O�l��S�1�u�J�>ȟL�ҏ*�����;_�G4�g�JN-FYdMj9I.k��Q:�1���5/�e�Y����tt�ٛ�K���� �,-Q��Nݡ�]���jS{cx=�T��V�?+��hq2d�׋9��b�^���h!�DX��03lȡ����������/�$U%>����v��Hk�@�nUɲ�<4)e���dͻb����WX�}ط;.�a���8��e���Ae�F(��|��E~0)Eh�Tk�K��������A�!����!m[m��'5Dj��]�0?3쏍e�%�-{��秨�]�Al���i�ZT�b�m��	N�y�+��9���Z�f2>%;C��ׄ�y�"�C��H� qϩ?*E��#<?��l=dǾ]�&����/��K��=�h&���{q���Y�|��S���./>]��UM�������x�~��hv�'��v6�19��"��Ϊ�PI�g�����q���~�y?����w��b1uU�Өݦ��/CВ7���'pP����r��m�ç����5�����{��L,��0k�F����cIT��$
�i�Y���Ɇ��};�K�L�ͣ�<iM��n]�ǔcy�����-I��57Oi�0��z�k`���~��T���0?jUWd�bU���Wo��r�@�4�����v���PA����9֫�iǚ�+����hG'�@�*N����g�êǈ+�Z��T���3�!E�6i��	�Mֶ%��rz�+�����:�b`-�a��`L��2u��kK�G�gt�h�v����z���;�����9�ZZ�Y�G�xS>@bx'J���B�{ �ޱĖ�F�u5h�;�{��W'��7�H��W�Y��"�Y�C͘�&B�YD�וb�E>��˦���Hﱎ���A�������o�sU`��N�O���E��gĉԙ��({�)��p�*�7!z$_��?�;�N
����s�a|9��V-V>��#-/��QK�� S.�^O�+av�.�4O����ӅLr����8��ɨe��:	!�$K��m��Ϸ��DU�XG����\�]�̏J}�3��: f��~_�#CH�a�Hυ����V=� �A�Z[�A�bB�`$QF�Ny+����fRt�-�3��/�4-,ws���t�h��YC7q�>�s_�f�R�O'�[D�2����z?EFߞ�]1���+;�)�G����M�@�#��j"�r��fS[�a�u	��|���f����Gb������E��u��,lj}ժ��b�6��odcC_�I����aE�*q�,޿�(B��W��H�%��6R�w^��;E�TlJk?y�"��2���nt[d-`���*�dE���c��<�,e����OrS�ժc��o���I��������ǡ������g���󡔯��"�%�A�s����:��}����u���ȟ��[�X3��������z{��8Φ�z��7a�!�1�����aW�Xǻ%�����jB"'���X��۪�d2Cj$�q���b#�i��ؽ��9ԑ{��t��?������Nq���~���d/Xt2�P���J�6ގ-P?��B�u�Z���5@���� ꖇ�W�m���5%6��� ��BŘ���R�S�'lY?�ZLTK���@F	�4y�2�I�Q������ح��%V����t�:x\�e6pD�U�<�h�������p������a�֠b�B�'I���b %k�'*v4׽�����I�Lh*�%b�7��0��G�����?¶�����~�^��K(~ ��ޙ.��˕s���yW��
�1�����oV��X���T�Tʄ��2�P�m��Z "��׃'���_E;�#|vQc閪���շ�`�\�ڿ�b��m�"���m`R�1������;hǀ���7KE���N�I,���Z|i�l!.��K:+l�C0W2Swl��k%�A��"�����}�1k�+5�,����<�t3$���u�;��OP��麔������5S����@�G*=�r�QPd<68RN�T��a'�A��{��|lJ��CL����t����k�k^�e�g"�{�.i�����ĵ�Mg��_�	6�|��Gq�/ݾ�R?�koP�50	�8�`|��5��VJR�%��k�:�'��m����AyR#]<���<�^��ҡ{��F�S�tK�}Q�k�T�@�]�$_�pK���Gk��,����t����j�b�5�v��7i�-��A��r�5�!#l%�a��Bd^B�.��A+?��a�v��� #�.Hl y��FJX$����Q�hc�Sx!G+�]x�FV�C� t6�G�O#F?5W�I�8@�㍐%���{�^e�(
?i�����=9���Wi>�}��ݫޑc�]}Lv1C��>�y��J`��
ϲ�a��{��n��Ca�;���I��QC�γNRB���e>F?�x�ĝ3(ǥ����1��ջ�N���r�BT��}.ɿ`�}Z�����B�<=�I��C�쬎O�ɇ 7��@ס5��{�&l��iҊ\ĦM�]� gG��|�ݛ_&ap4�[������T�x�UT�ä��!]�,��^s~�$�$x翓���h6(n��\@U�'6�씢�^�7 Um��n-��dsv`��\V_W�v������O��,t�ϸ$�|���~�*o���;)�N.��~����9��Pȿ�o�k��p5�c�r�"zG=xVH��|w�ީ�y&�,��У)k��e}��9o��Q8
4\\50�F���� �&��`�a$�7�@9E�m7��]#�,0�UW�+�]ģT������2���������]�_CH��B�e3+-�-�`�?���+Q#vū�>]���Up��oz��W��T�y�@v��Q9&+6<������:�3N�~�^O�Gk�*�2����)��oe6H�X[�cI�K��wn"~�lK�tS%�0�*�]T�o�X�Lm^̚����Wu��}�Ѿi�j)b]j"�r���� ��Lc�F��?H�`�������CA�lԫi��Mf=�o���X ��{Qm>9��Ϩs��x����e���L�eifU�����i��l-e%�L���x8�e����xZB;�^�EV�P�YSv�� y/��?-�(-7@��`a�K	��e����	1MTPC՞�fI���<Xp�t����<<sd_<MR=�8�>հ#^��+Xp��=z	�犰ű7�e�Lٓ���T��#-�m��7yu��ЇX�/`섻����USqM�B���*X;V��CE�����̅꩛
��)����
͎�~�3�G)1�������W 7.������'Ɗ�w�=��pR��d�.L�Nֶ�Ҁ�?�Q��K(\����D��'J��C���E���m����%��y�˸���^�9I��zﬞ[�/�����(2$��#�b��V ̬��������N�m�����E�B��~��U��'�5$��$��G�"{E��
�Pz2�����'�t�zG"���|*p;����f\�j���C�*Ԙ�V�@�$4sR�ڗ��7ǜ�<;n�����G�j�m���v��!���a��f�wd�R%I&ӳ�|,#�dWˀE�7_��_w��m���������擺ڟ �E9��A��aFQ�!Ǖ�)�j�a쥍 ^��wuK4ih�����ԥJ"��N���
Sv�.OJxQV����Ƞq
��/mnl�?�X���b��q<�f~��dM��ؚ�J�~)�M�f���;7A[�� [5{i�x���i���߂$,�0��⤎�S	*�Q��u����1p�R�ʴq�I��Zt3�fJ��_�2z������<�&�l��W��d%�6v�J�e�N���c�!���5��Z��߽��N�#PC���X���Ƀk�'�[a�+>���7�˗�-6��?�md����{�����iZ,��Y5�V�)��:�V��Qx��7���j�i��}t���!��M�7�*��(�ť�݈
�|vA)�t����h�vY
iO� �Q��odVͻ2�Zf�ʦR��ѣ/VeY�E#�Ut��|����'����zB�������A���j���ӭ������O��*��m[�RY�G�)����彽�}����κ��}Z9p�P5��?e���[�Ȃ<L��ױU�LSb�mJ��*,,ӷ��҂v���x��x�]Az������hzia�~z���R�5��?R��%���Tc	Z����_Ѕ���i
�|'��=J�V=c���5?�H�R�S��,m��\j��b�&���nJ��{�<H��j���ZA������<�o�v��$��6!����!�����O�r+�����]��4(ǣ%T���x�w/�h7v�T�)]^��x�{�zʋDʀt�i�?����0Zo �}�v0`��:�Q��	�����L��4щ	;7�v�$�$����>�^GjFJ�]��jrR<�������-���� �.�.�4mb�8G�nYɣK��Fq�g'�s�@��&>�G4	�{��UԶy_Tӿ�%2�˲�}c{���b��5\"�QAO {6�m~��]�����vg��D+��
�<S,O��ݲ&�c�3o�k쏄��3��<a�؊#Rx��T�lP���CuT'F2�� EU���M�ݦ��홻���$р~9=��u,}"���t��Y.�1UE�ɘr�e,�@�\�nU5a���^�&M�nY��d�]C��և���CDģ�y:w�>���=<�:��H����	$M+�m� ��$�M��\0���2�S}�:b��E%\r�a�������rk3à �J߳�5tp'rh�/�3v��/�< ���wT��*�\��[�:�#Pj�ǌ�U���e�"� ?7>3渙K	�|�Rm�/o)X���}{�{_ԏ)��q���g�� ��f�?���q�d5�z���u?�gp��t ��<~t�ӣ�<��[
�鵩5Ǐr�S�L��)cRp-����Kv�t�Q6����{/o\;Ȓ���c����4��3|��`�,�0�,x�m�|o8�F9��X�]�*"��4����=��5jD���� ������x[N���-�v��J�����bW�G������ev�㈫8?{|�~�3�z����yv���=��Θ;EEk�~	��;� A��i�'���cTl���-�+8aߛ~�V��E_%��&��mb�i�����E�:��0$�p������=ǐ9j��6p!N�b5����e�8��a��ȼ$_fO�%��������|��0/�{C|���
�`�Y[4X�Ar�����L�R��c[��w��@��J��ɨA_ב�-B���H����^���Rn��a��*��߈���;ٹ��aI\Ě��٣|��$ ��ƣ�.�Ov���<��|�/'�����TR-��K��]��-���Nx؛2�����_2�iҙ���x��p�
?��!M*�A���	O3��8�b��el�?#:�SŹ��F?G.lu�|4��V�Uݝ���F�7n}��2MG�܇����%f�����}.�A8]z�g+���"Q��^Y���';��	��>��è\#�.�g!�?�%9��Y���S\>�`�C� !�c-�ANV�����y���{sb�X_.�k��g�@$d�uQ�v
�|��$��O���V�k�������S^7��1�M�uIT*4�&|�\�Xݍb����?.Ja��6���L�-��LS�glUǠ�n��ςzp�v����|	�ye#F��Mr+���(C�y.�
YaYJ�+C�i��U!^�y��������)�O� L����g`�����q0��A ��d�敬Py�h<��1�����y�B���6���l�(��q���ő�"��"%v\������j�,f��U�Xљ�Z�hͤ4H/Aei%�56۩`�m�I<�扔l�H䣂獵������-��Hm���A���;�Eը��T���}�tO0��AiaU�{.��Aߏ���P��A,r�k�h$�u��N}Pa��<�ĕ�aAG��+�&G���B�kK�����T�ԣ;����?���h�vJ���]�� ဘ�:����h�\��vSK$��@U�bԺ~b�^ ��g�����*4�$��tQ��Yhs�:���S�e�]C��em6���MY�.����LG�o�x|�܋�`�>�l��������&Hg��[��Gc����߮���u_c��H�UZ
v�.3��ik��}pIz���a��B��������C}�D�\� �ch���q�w��[���kz<]7�t���>uAHp:klqj�^��V�/��!�녜�1:宥��y$�5l��F�-��Cx�N�w��8�Id�:?L]�p�GD^���f���K�q�G1p"g"�����l	����N��>��D��	x7���\�(�F�+:�^���U���$��x<[P	�������5<��"siVv9���Г"roDf����X��J�լZ�j�j?4��QH�G��C�vw�V�\k�ƽ�S���9+�_��==����b�����v=`�^T��C��ִ}r�\����Y?ar^�� 8��_���'�~���WlW�B�=cq�=�M���/�v��B~��7���7
��I��
Bb⟳U����wx�u J���b^��"F��vSR�Hg��:,0mgb�[s�8`��t�T��͢�`�-����
�Nًk��d��C�{Pa|oK��e�Ѩ*1�׫���
)�υ"�)�kC~�i_^x�7)��TTcf�-'�/@�� c��	-�+��6W`.�2d��"ZӲw���iW��{�����[D0\��(���c2�	n/��n3�A)0�ڌÆx�5\���Û�4��;���ͦF��� ���2VK��[?VD�YqP{��M��҄�p�^��ی��A!;�8�'Fr���e�w�k��c�j�UJ�-=H�v����b 0	�=W�6�T9�E��V�!�JD��,��������m��ߎyr��׏iw��8�J�q �UjM�
,j
�K�ٿ��T\ʧ��������6&mE�6��t�׵75��ˀ��O+�}�o�2�0�Y�CIW7�h3�VG��p�ʺ�}�E����r���\�G���*30�vG#��[^̿��uP
h����/��3�y�u����x�z�zK�����C�%��\����?!�jw'��¤��hbi(Yt2R�3����D�G����Ls��ܽ�lb�ā6��u��_�Iњ�HfB���]�5��B��prZ�����qv,�%/�(��]L�|�)!&���E~�6Ex2Wb�,ANfشV�;�,����w3�l��2������4�e(&�d/"�𲾟�%+&>��$O�)��E�v����|K�cןk��2>(,y��N�v���/�D5�Jn�7,�"�c�s����������^�Dq>Я��+�^-/�!�:c�G�~V�q&X`i�,c1G�� �fI7�oh�'��R�	'�U�a�w�-%K|c�����dHz�Y��A�W|��Z/�w&)���k�Xa+��l�����LP��_�\\����g�0��)��~sXZ�������Փ�+ܕ��#T�+�`�o�+�"��v���ge-�MC nSY�0I ��d��ev	2칧����%"�ޞ��o �������K &'7��=�Kqw25���n�dx$��2�ת�L���^�d+�d�`̡T���A�	��}�{6�I^L�2h��}�"�#~�o�r���ףۏ_��2>�T�vj<[֙����R����c����;��T=���Xs�v���_�e�D�l(�c�����'jVϝ���s?Pt/(�kN�Hgm�h��=����T��K箧�x=Z�x�t��R�3����m���Np�0��I�Jo �e~ܶ<o�ԝ����$�����	�3/C�tPSHB�V�!�5��6�n�/��'ﾠ����3E��w�X���&�M��|0�y�ba�'��T�J��քC�w7��:���C .D��mQ���lP�.0r�3�'5��Ѱa�J^-�>_T@��T
��*���?�d��d�=�q�:�rq�Q�\�yܜ�7ޱXà�B���쁜~'A����l�̚�
�T!c_D�\�7�*{ɀQ�Es�Q�;9��r���G���*u�4W˫i�z����{�j��k��/��M�L�Q���e�����^���#3��״ ��H~��#��X?7�+�(�*��v$w�B�0�x�P,��@���q���Kvy���~i�c�bH��A�A����ȥ�����&;ٌ�����V��;^�x�MS����9��1#
(K%�1��w�$Q-s��.��<-	[�?O������7�{~xϥ�V�P��(u�������U_�� �iW�)\Ѐ1���Ba�<���{�����\u�i�&X�ԊUJ�����C�̛��k��6tj' s���n�=SÁ5N��8���#�>�v6ם��m�oȥ�ȥ�!�[�h�C��+%*�v�?��O�{e�s/kV	RGwy����,:��V���,��%��N�n����h�� ,�ˎN%���6h���o����(�.�|t���?��F�����hkR>"R��ީ�� K��U��D�u���m-��V"6�����dHR��%t��j�A�O���N��[XwS~���@{M��}�g�#~��Y�X���77���/B���Ic>#i������=�S�q`q�E_�
��O8� �f��E���@�t�$��Z62=���>���/����H��u|��P�R�;{�H����"BH��n�Ƣ���X���c���|�Psѭ�B��C)=��sE���ė�p�K�Y�*W�}�/�S���C���i���K� Ҧ}1�g�[��A�d�i�F��57k�MM�����4���F �Řף��>��`N	g1O�g��zǧ�'�v��V#��L\ő/�ϴ�(����P֞2�q����-9fY��S��!�%~$.{A�1o�畇�P钿���-��u�p�	;s���tw�C� ����BT	HTL=k�֟�^}m�}v{������Z� ���vؗ�l2W��"�ױ`F�RR�Q^x#�w�u�nWh؏H�C��Kx�:����\g��J~�����y����3d̷xF�Ix��t�t��%~jR������Vv1�Χ*���"*x�A����`�;m}���2?K�ݏ�Ft���}f�]3�F��>�T�q&4y���w+9������Bة���`6<���5U7Ч�2�R�U5��Bo)	}e �?)�0M:�c`�����7�G~ױVc��X�����yRp�-��t@X]�a�"56RW���W�&���/0n���ڢ�}	M5y�B]{7 �:�����)e��u��{���Y�V��emP�:�@{%�5��
�'rl�mB2�_�D���Y����G�i),P?��=�+�ɩ��㭕`Z��(��IgI��' �Jvjoj'�}~<��y`U�8�T���E�+����G�7{ ��/&����c��Vn��p��.�j[iq<N>^FMC��,�5��C܎�cr���O�"��R�e�m �K �+5�ǂ�csA�-82�92M�y�����zo�)���)��
^$̚��x�/��8	���d=fC��բw�a������K�,N�n*����˻��塟:�7?_��a����tvs��Ew�\!�`C�>�pD�g�G�WQoj�(�y�m��C�"��Ȃ��|':lc��\��z'{�����	{�N��e�?+�F�%�AA�5O�XU9��^������ז���{�������1�����w�|�5۩}x�^�~�n�J2�� %4[_�+�����Ȉ[B�T�z���I|����P�4Y�B�5�W�sՀ6Vy���S� JX;�lj�'�$���b�vIDKQ�KF�NE��V7c�����	WJV�6L� �!A/�u[���|�O�/�r�Y �-3~9������^���D�s�lF{!� ��g���X�ظ�2��\�����,	��A�LU{��n�ϫ�
K w3ot�i�f?-��7"i�
�6Y_f~�:�kV��&f�\����<������	�����$Pؽo��������{eB��	?�H��m�nS#�R!�mp�a�ܭ�L�I.634��wi#5���-bZ�>�&�.}X�T��V[�T(���'ri�m�s�p�уe�e����"G'�(��-�GR��?*n���?57Z��BjI��\�rߓ��x��d���'b5��Xh�SX������cl�Cpw���U�����Pm�t������x������{� J�1��g�r��γx�j�i4�3�k+'�����`q��z�!!��9L�Yl���_6�do~^�s4�\bP�7�p�6���i>��"2:6�����:�0�՝�ɻ�� c�+1���\E��+��<���:Z��X�O�L�?&2�5<��A���=��o��#���GA��C����U��,Ep��u�r�WL�uN��{�u-5HԠ�M#�TЁ��-� ;������Z�
%�����Bq@��Y��O�(	�2�ϵ4�]y"3��fnR!�C���F��ؠ��: ƍ9M87%'�����nj��*u|�a���`/n2�u��]�m�OÀ���R��/�į���� V��3e�(���0�����=1�w�b��n�e �]ل��7���R�L�5��t!+C9�;�'m{�XN��4�M��srl����$»¡leⴠ�n��5D�,�LMr^�v�KK�I�1�_�2ƴ=p. ϛ�*���ta�ӭ����d>zn�T��qb>ް�:>گ%�BW������(�=��/�y�Rg�/�\�@Ny�;����A�p7v}�xn؞��4��;��f;���v+6I�?Y���##���z<j�}�Ī3�.��_%G�]�� K�����U�g���腅(���M�L'������'�]�!K�9h���#!�}1f����o�o}*!�������|�Q�L�C�L��k� ��UJ�����\� �֬[6COP�#x�q��ou��4|�{v4�CȺ
�d)%R����Њ�h���ö�*���z>1����}wR�kT�1�vqW�H�r>p�������Ą>s@���3Z�%-8`��+���]������G.Ax�F1��j� l�&\�sT��>��V>�������`�����89������$U���bvc*桗�IT�XR���(����j�֋�S�1���9.�?e䚷�bO����P��٠Rh=�!�L���/T�np�;��@�r��� |��V��y�U1�]���_�a8�	wh���ի�yU�]~����8��&�n��2����<M��h�$�I��3�5�H���VA?n����3t���ѐ-M���n7��G)-�,������m���Toc�"T!�arT��sst@7Rm���`�>�H�?�Ű�nѥ�J��$��ã��	��; kTp\��AR��N`f��
���+ۓ��;��K>��>�oo�n�=6'���v���l��ط������\.��dޗu�Tâ~������u�鏩!�;��[b�­f%:��(Д���j�I�}0a�'?
?���q�y��w�'�
� f��ktq�S�p���𦼾^�_^�(�݆3�����?�&"�(��j%�s�xN���0�%�W��/NWA2��I��V|/�O������PyN��YK��og��]f���"4e��u�]B�O8�����Y>�Wʙ��(�I���$A'��0���v�`�q"c�_���ҩ� ٰD������Zij�3��R]���J"�i�MY����1���"���s��a�;�M�$*�#`�>%?��m�깨�;p컕����ydN�[�	y��.4o>֌)>\O�ʝ�+��b�
�a��;eܖ�@�d�>�p���D���]�ն�J��D�
�.Ą���"����3,�����`�g_gak��nl*	{�o�W���Ts�F	oBO���q{�l��V�o�2덳"���"�{�'�������Ʊ ��Iv���K�~|�:Lg�s�.�柸x6�ħ�M��
��1	_kW��тDV��ݫ �G�v>r5�׃4�e��l	o�#蛢B�X]�"��=�t��[=<�slE��g\fPY�ށ�G���5:���h?�k��<�:�^?�k�:�q��F���Ū���c��{�m �οYXj)�ҿə-O�ꠞ����yi��s�$��m|�
���7��:��K��7��N/k����A�j�Ɋ����k��%��c�^i{�4i��7����2҄���:���`�r���c��%� ܅*�י�:�'���8�}�;Z�	�&4,(�cf�5d��ܼ,�x~������鲣	�E�dM��|)��Q���:&T ��f�%~ht�JO��+��n�X��V8H"'��=�&�̆.sN�gSrqJ�*�%��3�,�C ka��qsfjd.
�B��������'1CZ��/u�Q/[҅�#X� �4�<�$���<�����'w�C�������VW<Fx�1��l�Q�g�)���!��Ls�"�hB��ze[<�n~CZ��,	\5��׾�#\֒�ܪk�
:1���'���n8YÃ�X`8 ����	÷����o�0�����N��
z ����$�Ձ\ܽ����:#�E�*�>F�� v��f0�9��NijK�r�S�<��[�4	~s#U>GH�������xe�`Au�,��'�

_����cl����[��
�\[}�V}ki� ?!��{�*<�Vt�y��o��
'3j`��z#�*�����/��h�;�R$���R��ꝳ��+H�<���*l=��E	�r���~i������1���;�wb3����e��7|K�k��R��DC�qZ܇��yb�o�Ξv�����m�٥��!�7!aJ��o���Ep�2}]��olBs-��6����"�e����?��fi�4��z`t�KO�i�C��RR�� �q��Pɔ&)�{w���Qq�=���[{>�H��Q5Pڛ��oz{�B����Ո�3�һ�G�q� �&zW;���[h�s��9�#���R{8J�k�,O�$Ҥҁ���-�GE��=�*K�t�4L��nu����=�/)����`���G�禍$��B=�A6#�����.�8B����=��'���$.�5��j�1�  Ku��icx%�ex��;�Ƌt���z��UB���y��ۻ�7iB�A�+����+����ة���J#�����+�q�^<O)y��\i젹�6���5�����;��\n�d6ʧ�7i��Os��h��6J��Ӈ��4�\	=Թ���s�OE������+��)j�\*X�	hM�O!�+�H���[�q���Q�`Eg0jL��ڗ^XrF;���W��B>�?7^�����mĨ6 n�m������i�C�f���֓��D�R�Oԃ�<S���ʰ���ȍ����(��K=��P���<�3��x�N���rE���|��)]j���ڿ���XwE*�Z�'�w>��pG�vS-�Z�nr�B�~@�S�}"5����n
���� C���뵎�fT�>�m�X���Y�PfśwM��;7�09b�R/��-�	�bF��裿�8p�ţx錵S��9�*r�/iﷸ�q$�	L�d��!���iY���ӧO�l%(Z�ΰ��ש��zc��w���7Dy�e��'I�֝��IewT�$�e�0�X]�
@�A��.I�	�ĭ�w�������.��|����8����r���Ӎ@*�!�� �ɉ�%��zJƣ�����^���[�T�T(G&�����-���:�um	�h��wER���A��i�����
'1���Bk��B0�k-u-D �����v�[��ϭƵ<�/�	����K�N8���G�Z�q�J44ж��{ ��Uz甥��e��b6� Lh���$�벫	^��A��f�?�*^sѸ�9(N����D1^��Zޅ@��'�)I�F�7a�oϥ/���s~S�C��Om(��āi٥ɥ͹`���4�c{Jg���ev�G͉��Y����������C�k��~��Yl<JQ�<N�vh��m�����O������E?)��������"���p[�a�\N�*G@m���^A/��F�J4��LY^DD/��%1e�Ӥ����A	<�r�o�ݛ������ThA����q��޽���7�hDJ�p�v��P��0(�E�T�RWr*(�������񊠹ʀ�kA#���oZ��E-�!��^u�B���o��2�l�?��ӄ����ns�-��o͢	�M�U>/�:��~%�V�������r�X����+k�(02��ճ��o���"�� �h����͔{��gQ��������z����h'Z`)�O�n*p*������r���;��װ� ��A���8� �^��Y�S�)����J���`���Q�ԕ�>b��r�4��/�{��B��W�E<-��&�K�Q�Q�[	�*�֛��n.��m�*ʆm�pT��xMݦ�IK�E�J��:�=�z�09T%�2c2������<��9��\4]�P�J�n:u9��R�������rO
JI~@�ѻ�d�c��"�A�\�FEgc'_4��" �[�P�ą.��k�M�.����/�����M��yu�q��#�G�|
��}i������[������7�2P�q�<����z^�g�lB�y��=�䐡�
z�6�)��z���@K�hK:�$s�,���c L�
':ph�F>��D�-)ϧ�J�i��xq1�d�O ���>��xU�C�N&ua�u�o��9�!u��j+�'�0U�a����p
��)���:L�>��@n���V��U��śf����"��\r���m����6��B�"�X޻6X����f뺬���f2���F��Z�7�z�ɇ��{��>��-*Cfv����l�/����Q�K(c�ppW�L%��I�jӝG�e���D�[(�M��[�*�r����T�=n�g��W�A"��Zȶ���R�0@+w9U/�&�P��̲�ԋW}Q��})b��Fj�r�3���E�-������wU��HE��0�e� �O�V���@u��o2�m���o�����~I�q�/x�U��ąc
�ҡ��sA%��j;�&)��=Ia'��c���(wf�ER�,Ǥ5��v�Kc�K ����v��f�t��8](�^���u8�rw�Y�f=��(eY�ٔ�c�H�^zRJ���m�%Y�Y�R�P��Y�bJUx��|���7y1�F)(�IR�P��5��N֣����
{�w���)�H�&�!�XDr��[����3z�C �����eT�r ��m�����M�� ��f<�$9��"��pT1Pl���ykf(���6�LC�g��C1q��֠F|:�vO���+50�Lڛ+L���G�	c<�G4����|�
;�'�̀�m��6r���2uBt�#7�^B
i�]�G��+[����As�I|�Ni1�}�mS��@\�L/.�Uz�[f�_��M=�mb+l'x�S��|r��� 
����z>��f����2"8�9:��(����\�~}����e~�B$3�B2���ϔG��\�^�oU|�͋#^f�x$�ݧ�G���:g��*�>Ȏ�M�0�W����S������2-2�_�v#}�骗��ND���5�$}�'7����)5�����44�[C������A¾�v廤�u�2��j��˟���kG�s��l�.��gx�{�Ps#��Q��k�q�ix�jգ��-ۘ٥��,޹��3���f-Om�N�p�����-ɇF�p�������� l##��;���L��L���e��;������F]���2R J�Iu؛���_qlP���G��o� mQ����V��z�����̻F�Y��/Ai�QL]	��0��c!����,��|��`j�Kh�%]�2|��'k8�^�.�O����a����w�	ۉEe�YN �R���JtP�8�<:F�J�ޠ/��� tT�oQzG����\h���H@y>��p�w�UZ��{_d�-8�y�8�9o7�w��ǀ��^�xR`�7b'��}�UtB�"ܛ=P�oŭ����B�-�h��YԻ��Y`&��[U`C��ID��(�����L��[��0Ø���" �S�����ȴ���O:�.E2w�	\�ɣ� �4�ZS��x�\�=x�/���ESi`�oh������^@0?t��*9n0���D3Pif~�e��8���$0��[n8��DT�O���.s }֥��x��_��4-�� ��H�W�2P����� M��{͇a Y3h-������h����~\L[��g/a��R��b�d�q Iz��`��z�Ml�Wo@W�c������+�<�'# �U��uL�vG8�̳�Iٹ1(&��:�rP������Wc���,�h���}�j>�a�ԭuн����pQ�B�mˎ�a?��p6�2/������Bg�ÿ��ST�uɜH�[S��
H%��T��������N��*"?��7���ё\�@j_N���Ir��('��)x�K�N^�;I,��n�\K`��.���^���*T���ZSA���n]�/AZ[��Q�������OG=�hg����9Kq��섻���%*�1`9�Q��(?RP9G�y,E������; @(�`O�~��� ���6�]f�U{��N��C�$�92}��p!|��F� ����7�N���N����Z�:���N�fO�����U�X:T�ǎ0�'�b�Vd��:ut��6QGh. �+�>�}!�<��/
i�?���m���$�!�U�R�e0B�&o�+��)A��T�*�P"��qo��o����aS���g�a��1�2�ؐ2���~�kP�y6a�R�-H+M��R�-[	�|V�;Gt�.U&�A�8a4���l�#sξ����q=��[f�
�Y��z8��|�/���^t<�z��|�L�vt�J?�5O�B�ϣ�r�5Vֹ�gy�h &�f����l ;{w4{'n��S���dH,�#�I�ֱ�M� �B��~Q���;?
-_���� ����'SZj���̡a�׌��Ax1���j~剫��h�,�c�������b� �oT�pE���,ah�i��n����'���C�k1Q����}�~S0��3g�@��ô�/�/���:v�Y�'�Uphdھ��ꂣ�m�ؙY���!Y/��y�W6q�Y�����.ￃ�攠���x$q�~ݞV7�#�x� 7�pE�
�HIѲ��c���%/�����U쥰գq��T�q7��zE�>$4�r���ٖj��)K��E�$�At-�\�o6��R⡘��]��aW��He����mQ~q`a�$d��ym��չ��2�PxT��4�'	�⿻m�Z��1��*��ld�W��3�g��V}X��@�hԳlJ~���<`�'��UwFݞ�ۢ�IR��Ђ@ (,����;�,�M�$���C�ӔT����P1Y8,t����=:S:\Ⱦ݅�t?�}(A��C&>^�^�� �
�i> ���� Q�N�Cd7�fIn�(����� �e���j&�^U��ӏ>L�%IQ��^���~���V*QP���Ae���ީ־u�ʅ�`3:��;O.D3�*;\y��ֵ�}��$Θ����|�~��w1�F	g�]!|�hu){z�Ӿ1�k�`��a���̃λL�WB T,K��b}J��8�!x�s�ꨭ����U���'�Ў�'TW���P�A�:�b�<|�_R�g��"A
ё����b �:��t_�5�hx���t����b���œr�DO�MEw�I�Q���[,���Rv���og�o��T�-�NѾ�ɼ��iI�������y%RP��ъ�J?Y�� /9�:Ap�����k&����Lc��&㘌础Y�0��bT�KT}+��b��`Zƌ�����³�P����C�X.3�\K<5��� Ԧ3�J]Pަ�>O[S�?V������B�P����ho�w�F��q�T�3��7��-������0C���>B��u���9�
J�}P&�>iz���p����%��FP{ty)���a���an��sJ��dߙ6Em��-:x����L��f\%�R��l`	�~=��ar���'Ԫz����Y�(��-MBh��>������N�m�S�����N[-�CmM���a�<\!6��X��Ta��3��@��#�b/��f����3?��������n�C��G��EFSǏ�Ă'`X[G�`���G�j���k�f�]�7�q���.��~��Ú���A$M�V-�"���5��//6(�"8��w:���KB ,3���1%�܀��L�}�J��D���>���sC�Z��?ىs����(�Q�g#��i�b�ihة�l&!l�q"!�����~ek;>�;ɣ|P7��u�^Px�z(F}��`y�mo�ᴋ��/;@�M}Y�����/>cE˶���C{�B|�cb)g4)3��nZ-��3�T!
R�P�HyK��<A{�B5,@�
����1TaHO�}u��l���q�y���	.`X��[y�����7JOC�UU��Qk1�����|s�OI*�	�A��J�XDv O�&���j��N�i`&�����8(����a7Mbs�v������K��&�n'�^�@��ـ[���$j
��:UK�_��P l�p3*���D�do���l^�|��	�|��k� �wwT	_���Lٱ�A�ODZ��d~�{[P�+�y|X�V���>�P�Z�h�])z������ѧ�WJ?h�?S��󭝢D�q !5
|��pe�^�]]]*N�
��V�H���r�P�&����N��y\��,���|c����N�	*�m���'|n�,"{=&)9Q4����$'f0	�_,T�D�f�X7G�?r�FvN^�E��YP�[f��!�W_�]˰� '�۪�FD��M=߸w$U�}�2�sfI�Gq�)J ���>A���j۪j4ⱒ_7ڦ���#>:Y�� 	�腙ڎ{ڪ�Ɨ�G�ˋ���ؖel:ɒ2�>_�ܚ�E��|y:�"��Y��(W�P��J'�^`��4.{=�[�J����H^|񗐙��qJ�� 2�6OՀ�FM-���;��J<e�΢5�áe�u���y��1U�̵��`ָ���;����U�-���o�;���͟Nѡ�:O���GA�z�R#;E�NZؕ���ߒicω�s� w���5@�υ+U\�g?���p�}_�A�|�,'�,�N��YR���ק&�� X�_`/���j����Ɲ>ݕ�����y�.���1����I��l*{��<�%�ψ�BӘ</�NݖBĮ���W[1RL���H��Z�u�������<$���[�Q\�Y7�\�B��on�{&�y`�	��l���g�ԫ�\�ơ8��h�C3�Ղ:��pXD�,i�P�}yf,����`ؖ������ [�ة����~�SlN�)#���4f�]�U���!z�X}1�(���3a�L��ط�l
�*�������Z�B$L��FU������,IM�8�Mv��^��S:��v/Τ��@_���U�J=�;�aL�e��x�p[�@\�Ey?�a�����{�5~��;\�=�w�PQ�)�4I$��6�j~�o"�y��������\����0�E7�S:�����^Y�+.����RW"�"B^zB�� ���$�)���S��GA���{����V���:���O$I������B19tdU�?��\wP*�DghCxz����y^)�ٻ{(�o�S������9�ej���a�	�{Շ�Ǉ	��s��p�Edv��4$��H�'%u]�Ǆo�2W�K_��B�\�\��Η�;��NRg��r� Q��]��ݯ��Su��OL�?�D�e�x��֣��'��h��?I &�t�r�o.��������
�Sk6E��*]و����b�x�-8���B�-g4����β�LlG�7�AZ:��P������ b@�"_Q岧*���QAȁ	AXEp�I�����~�rF'kʎ��Q��u�Dǹ�g�u�bw�����\�D�!v���-g�H�|�J>.��}]�6�K� �d���nl����P�I��l|����g&�ޏfG�]._��̥6]�yq*��u�uw�\���o�Vx��]��ʟOE�����*�E�R\V�&�Q�ZIZ���}��1	+���Jc&�&�����v�g�d�o� :�0к�	Y>{C>/�
�)*J�`P1�*jV�C򹇓u�
���?����dbP;:{˱ޓ`3J��с�!���$U	��3��)�Mnf�<�,]H��1o�-�Z���Q�l�Fm�bخ�D � t>9�G��'c�e��Kc��B���!7���,�)�ȤK�V���]�s��Z/���u��Ug�y`ًO��.-�-��L`=�:��|b���H}b7���ʩ;� �r�1�,�,��ó]��KKf5�*����ASa8ót�~����!`���l��ԁO�z��M�~�D�+l�[$�^D�2�-��,� ��zc�����>�6��ph�p��JNc	�`*F��2"T�kcd�T(v�A��A��7=ua���en]&�,���vq|�2^�U�ы��Gkr{�B�aA�n���D�QQ��PޱDn��{>���~n�p���J��"���{ç2���BL��
�WZ��sJm��w���$���=�8�kE��هm�6�"Г��*�C3�ޘM6�,���NU��s��7'c��3(�U�f�4'���欲8�WC�zD��L��\�ORI�0u���>��ۅKR��}�,rw��ͣ�H�`E��BD�MW}o��FE����ǨC�G��wc�'�!Ioj,��s.��g���v*t��d��&Q�g���n
�J�R��NMb%z���-��L=#��\V�g��l�_1��?x2��y���a��8��������߲^�lze���y��5SF{��gJ�&�{hP�G�dg�#��l����#D�:�*����Qk�G�I��E��|�SG�2�`�$���J&�El��ސ���A~�)NƘ�˦�j������e�C����b���6�����:��G�>��O����*/e�!fWW��V�]�o��z�qMS�����D1��&����+��
�h���"���̂�*�>Z�d�1E��W���N�� �[�䅜���{pTQ����K�C0��1�O����������X�����'y����_�b휷��9N��ƌdXq:H��f�>K����:����:S�i#d)����`S�q�ک'q���S�,�Or%�[$�&{S∔�~^�b`ȋU�1�[�n9B��e���srS�rB>_���|���*�|��G&���R&��&n}d�۵ &���C
�:�^�
��QJ�4�{�/��#��ByYx�g)G�����D�-_�����Y�����	�^����k �0��ɒ�k{am�|lq�zz�"Vʛ�����忾�{���F��Ф�6C�ts=��#<������Ƞ D�(Fn$��KrB�H���hA����w��)�EjEE7ˣ�kJ�6d+�(�#�X�)��.��n�:V-��2���w7@�"�PN!�y�_({93�����ͳ�����A8�"�ݐ�ḻ2gNSv�b�M$�Џ������"��pq��6}?S��:!l؃�݉9[���l#�~j`Y�Z��T��ȸ��&�3��$�8v��tS�y���L�� �-�H�y�n�\�ҞK8��A�7�y��s�a��P1��%�db��\+�x��,iл�b�&������ʔA�u�:�f�;��§ߋ[��W��7���5��o^���Qg��&
���p��s���ؗ7�|#,"��[%]�|�"���ȫ��I�H�y�����ބ����z��n����T��)�Ո}F`��.���a6�]�d�X�Γ�>㝈�sqY�H��?�T��$��Lzg��/O;�
	�a���_a��g���}��:��W�n7����ĺf�cO?�k�KA����v76*z���)��ZJ鱲�XzoO3\$Z�]5��'�!��	���:�{q��L �[���b�D�B�d`�-��x���]�׫;!�[�̡�L\�5~Dy��bŀO�aF|�����lݞWn���jH��؅�5-u�7��-��x��b�V��r�ܧ�-*Ŕ�V&w��<�y�/���8���l>|]��Tz�i2ت[�J�R�ӪB�_���CP���¤���W��"� �Hi�F���~����*q�ߠ:��d]�w:�s��55�#@�`5pv\���(lx%��c��>����>T���f��Sb��{#�%Ն�]�UM�s�ډ���[sW�O�-&#|V�Uߝ2�3�M%�â������l@�>�?�?�į����jJ{��t��������[�)�<�l���l��E63N/t�;�?�uT��O��<�x��Ҧo�j�LL��j��ԩxi���~�n����	��N��!U��t��D��E쁛���ec.��Fh�'��V�ӹV|�
l��h�p!H�;Mؿb���P��������{�9��H�|�j�]gf^�kY���j�MΞ��U?�ԉcCL����X#�7��4�;�m�6C�c���� ���J�3/ħ5U���p5��Ş�
�Xo�G�,C�Y����_�4h/z@�S��bq}������"@bx�e��7�����|n�M�݄��R;؉�=������#�̓]����4x�ܰm+�C��w��^�U=���E�g!,mG3�WǕo��Trd/o��p�
p9Ҟ�T����R{�?��<�ԗ;�ݶ� �i����5 }�Dۄ���7���e���Ur_���Tu6`kx�d�_[�� W;�G���|�	ӗ�������iο�?�t��}���M�q�rm\�v새D�9-w�%�Tǋ�~02l���A"�5Xki�3N��ba^�4٢<��7�~ѡ�.�J#�������F�*�lU�S���ٞ�����x����E�7�W&��q��]���-f�U��8��oCި�McX��K��D�D��~/��x�m�m�����ȠJ	X͈w��ԍ�c̓�/�F�PPF��6/�x�H
��/���ߌ�3��#���F����W0+�Α�
���(
���0� ^|�q>�j�@*^�C1% ������V봳=!Z}
h'��s0�]_�&��x��Օ#���^�2e����9�N��������~��pG~JdL\pGр�cC�U�	KkA��,}�=M��8;���҉s��Y-��
���`R}��i��ART��\�&���q��Ѝ��f�$�vH:�<�5�w��P�y��������}^տiۨX1>��1h��y\o�����*]��3G��2��/��V�4x릺ka/�ݡɆ���&�/�P��B�f��_ JKƅ1�ʤU�����+������ڝ۩|}ͭ[�� �Z7Y���4�������߂H��v%�'��' 
}� iy��6܈�����r�FE����%!�M������<f��ܝ�tb{V� �V�О�1���k����/���T��͓l��� ؜tI��u�V6�O���i>G�EvKp��p��Nv�-\��V���ǧ�O�{{�)#>4;Bd(�v��]cЦ�j���WGFTP�ez��2~I�[��-��q�_�?s ��*��L���jY�D9���S��ViӇNhy�so�y=�tt�0"4-���j�v���.����Eq��QYg�*Ur�ҁ�*xCj����Fo�F�[ ]	�dL�	���v8nl��xI��%��jz��H\���{0�A�S�:H��|�
}���ٴ�D.Tcdz� �(DS���ˣ6C��
;��"�[z6%ލ@�%A�gw#N�TR����'�v �����c�d/��'p��оHĴ?�|قX�)���؈��m�_��5 a�����li�/�k"%��f���ƺ�s��ʖ���y��fH��c`��\��4�g�]��g��!uD�Ј �}���z�����h���s]�
./H~ƬP�d�dE��e��Hj�k��/4����5�2"+��۸6a5��+=ϻ?3�D 
��њeg�
o�Td>� A����,�vӉw+�^�,������s�b��~����llX�&λqE�h�-��@�w�Va8=�hZp[������[�:y�b�L	~��p�['���f"��5�JĴL�F 	��Ԕ�~�Q�l�-њ����[%<)Lt�^��i,�(���ȡҡa6����[o������瑪��31G.�xA!��އa���'��B,�m�W�Ȧ�c���tI�p���ҟT����uMv4N7�� 
C�Tv<Oai�9�F�V`��P�*#�\�@��W��J����4�>�a�L�u�/<`�؟Q.(�uYR�
x9��O�]Z�l5����Cǂ�J��O �rGE���d)�-��o��x�m�`udF��gC,]Ή��GT�ɾ�s��^��'C��ʘhV�<Ԕ��q�W/S�$0O~� ������4����ۺt�5:ԕ�UD��*���1	�9$U�h�y��fN^�)l�t�����>�vd�'l$�,t�\��HR捀#K��?�5�~|#z��n��sl�@O���b���ۥ}Z��Gt�d��H�Ls���q1�\&^��K.X�(�mEom��F�u�:
_�䢍GK����N�:�%�L�]���k�cZ�XH&Yi������� �F������e�>�؍0���ߌ�b����5v%_L�g��4�s����`[{��iD���w��TLQ�1b ��Kbs̀1���2�	�w+��$w��C0�6�E;�������U���i �a^�Iɉ�U�����僃��2��}�����잘��KCL �>So?��"��'��k�Ľ  �D�K5�(0^���6�=�W��P ��o[w��iyT��,i᥺{����1
Y
ž�~��ŝm��;"�i��^��{��r���T�{�.�a�[T�X���Z)��l��ؑm��1A@^�*aCO
�0��T87I�:�����"������l�C4]:��d��1j@d��b�CA���c��8= [�o{�x�l	K#��aAx������X#�i��������^�+���E�/�����F`�����sOM(��H5Ƌ�r���<��$�h������p��C�g�ӊZ��M��V�,�1��4�j�jx��.�x}�-\��x�T.v+"���hbv�i��}�Bb�;�r�
�Fw��)sG��0o�	m�t�֑���?��&u�(����߉�]kV�u�ЗV��.J\^-�V,��Ӡ��V�*�W�|d�K�͏Yu�8�σ��7tRvrw�BN�]�!	w,�䍳M�܂-�?"��8w��*�nt�L'"�S�TP�3�J�߆+9#�Rn�֔[� ��;�.�*s��Yw�ݤ�,�+�[x�X۷���6���2.��Ȫ�S��jE]~G.P����t
�S�i�"��^��Q�n�ʣ���+)�r:,���wS�*��$^+*>c�]�{A�ʟ�ۡ�^h��xj�K�e�wm�h=�R�L���ˀv
��k���J��d��̎��lD�~�'^}9?�p��04==�Ӄ.sf�8��l�+����ic%�BE3��Q�DB���=�؟�I�VP�;&5��h��i��/z�NA�(�b�u9���1�T��V�`�c���4�N�K ��)nn�}S7����hW�ǭ�Ɯ�6l?!Nƈ�s���(6���p��]��b�e�N������\�	��X5~�ΐ(z�C�{M���	�{m,E�ݬ�#��rS���:)��e꣧�t���횶p������r�a��lˣ�@��ѽW��T0�L��G�Le64�]Ǒ�o�z�m�7=��v���L�8�[������ �]�yq�.�$[ֈ,���(���˂��e-����f������d֍�&�콻��l;�O�,������U!G0�����NQ���b��Y���?��
�Z�t�kf7wfs�K_�!i�Z��#�,�;����yc{�zw�{x��c�c���I�]S�X8hn9�����5�bI�
)&Y3W%M��Jbo?���u9�o��vh��j�Zђ=؝����D�����Q`A�>��K��вHK �\��+/5H³�(:,�tm�62M��@9�NE��#��?�p:l����hy�d_S�`0�����D�fl2��\/�?�AwA��������O,�d�x�ϲb��D�gP�-��<�AeF����zo�ٜc�,6�zƞ��`H�3�Jÿ������,>���ͩ܎�QA��_�N�D����z�%?(#MM$WkJۜwJʔa`�*�&s3m��=H�Y������N` ���W`�ңoF|V?.�>��H��Q"� (р��e�r��Ʃ{�+��8ʓ�h\��;B�E�J��j��� ,��V-t}Td�!h��̿+΅=E��/��R7�L=J���I��%8�TðC��m�lz�Z	`X=��1��*D_�� ��	����n��T�D��Z03u`dR�ޘ
mv���ϳ 3�x�_�4�|��Y}�ԃ��e�oc���q��K�'�T-�\w�Ή�}˧��Np������)^Xw?���ja鬆m�Xҭ ��y&`額ٖqp�v�ݴ����o���Y�c�vb��>g-˵�@#՜��0E�|�hDS��d0~�H�hD�t�5w	���5�7��뻘�b�f,{�q�A��)F�HW3y�6�I2
�E17�"��|�6�#5:���kyԺ����3[�3S-��ݚ�=�^����c�l���Y4��s~eq��؉i�5��j8D�jD�b�w-��A�6�p��&p-�^pW�s{�4�U��f��I�7�1v�m������kr��fwyx��]�`�Y�m���we�J�E�yT�?O��m�i�t�� 57��|��8��%�He�>j-o�W�����b�O��m��Ej\H,�u\�j��VƝ/��\Tfȭ]��2Ue�[�|���#�mg��_Z�5����]��N_��_����f2UR"����NV�A�3(*0ɱb�`�6��H$p� � �^��3��m�S�DJ�c*E��ϳ��T1G*�I{�z���-$�&?�ǋ�=�Tl�S��Dϐ@���)+�]6;"\���Z��5��!�j$��v-�/�6�K��Ŋ���a��A:�L�<ӛdZ(r���ͩ�U����M�����A�U1O��>96Jh��>��H����EF�MYRz��f���ʄf��A�k�I���|�����m('	@	��� �O����q�ћ���}!H��Ml�x��&���Y�u�"���O�}we���|���1c�l�})v��H)삮�\3���mv%�y��~���u}�'��HYy*�-1��܊*%6��\ZeXv��	v��jy�|�*I�o��x�$��ʖ�����7��a�mK �Q���ߖ������q�j޲�/H����P�t,D��H	?X�Q���n��y�6�vnl�٬�D�j���,��箧-t��&&Ëm�H
�? #�m��և�t�ְ_C����HM�s�©x�Ѳp͕X����C��`0���W��6{�������'��t��`��Y� t��րp�S	|j�~�`��eƖ�q�pA?��~��=��G4ۿ�&I�ei?ѵc�-š1�aQ-��F'����&�&�X�x��~��(5����Y��rƶ�<i�ȾMՠϼ4V��7�+�73� .���y�II�����~�X�pt�NYQW�̓�ي��{)�<U#�2.�O�&���_n����0:�a.I�+�6�Itgm$�k���x��~�>5s��[�.�0�ɤ
���4�y��߳������ם�d��>�+�k�A��)D�����\nG��	<�^�"@��u�ާmS�#C�tL�K�F?:���2wA���t��3�b�%}�<;+��O:��*��B�?i��v��z�Ig!Y���������)_U�CV��K�� !��k��~��/gdvi-��c�}���4S::V�93]]���Yɂ`��j���w�6݊m��V�-=oش.���ı��(P�P]Ւ��j��M7����#��6� YG�dD� �B��%��sЋ� �_������@� pl�m�[�N۩_7u�3�ZpE\ �$#C;��d��0:��'�j7�8�Um��{{�+��L�N�::V���5���,�pΩ��Z���O8��n��=��ݩ1���ߪ��H���J�0z�l��4F���G@��+�{�EVb���D�ϵ��������O�P=gl��+��ˮ�U���s(�y�9c!"�&��O�6yx����.�I��?��i��q�E�@ڒ�<x�~ooG�b 4o���]O�X���V���7gv����$�1���m��A@A_��8���+��t��:6����mGI�{Dw�KL�3�t�]˟���'�"���`����|�v�y��E�O�ac�Ua���Eh<�6D�9)O�P@	O����{T��Aeх9.Z���D��wd��g�܋Ġ��/)-W�M�t�D�?>J:��N��[���&��+�4C� 
��1�1�<-Q/ ���vyUI�]]I&��]X�ǉ�b2�Z��4k���s����� �kǄ!W�t�5�&�[��W0��"K������0D��@>)�``�(�����r��<j7�M��R�Nj��C}2�U�w�\�
6�;P�x6�R���vdW�����+#�$-�'M���˴]�����۝��o�MYXF1�����5����H�d1�~�9��{q������Dʲ�z��X���S� �5������כ7�SP���c:޶�Ӳ�` bO/��������OߗA��M�N�"ڀO-��h�@|���Z����,Pj!�}_����X�Q��nc~�it��7�Bvø����yؑD�7r����;�
{��Tv�������o�ϴ&�V�#X��J�>�82�ٸ��G���3+j'//�ƴ��P 	�7x�L�&#jO0U�ϸ�f�:T�U�b�G�k�;�V�4˗	z��H%&Wʒ�{�N����P�}�n�7�@��U�!���}�q	�j�&��!��������Ll �c8j���ޯң�nl�FN�a�H�.v�F"���߄}s�W�U�pkdV�?b�1_�� 	�2���	&��FI{�;6��M/�ԙ��T�%n���յ�D���xKMvarE�Os��pU�k��c�u���ޏ��t+W��@�Ɣ�� "�lR2T�	���'O�!�_x'�ڡ�J3r�H�@9z��O��>���:�û_�W̮�)O2.뭒�``����c�X�]�����,��ְ�HI����GU%��O,�#l&���C�V�K԰Gq9`�E�v&�㙨A.zy(�������D믵*��&��L�V��As��-���n4��X^[ͺ��<�*�����{��Z�b!��d�7�����(�t���U͐i$�C ؿCa��kg�%!�K����v�[Ԣ83$r)�y�xL��VX���%LgI6��) �ӳ2j;%@�o@�
���"�YerŃK,�_4�N�,)ޞ�����+�͵T���@����~`d��\;������%���BC����7{�7i�U϶`�U���4A)=�α^&@`P���y�1*ط����a���(�?���%��.y�3^�h(/��Gm����1c"q��w��<O�A�/~�F�bc����7S�R��rD�e��2�P����r��{��x-���ha㻲������G�C|�_�" E;�FHh�ha�$C�d�CE�N�l��N�Z���`t�)(��Ac�	'��(ZT.]<z�/�Ҫ	�io�S%�h��u
�>���U��+���ԩO2g�c��D�(br��Ta�r�PӰAں4�s�0~�f��~�GX�;�`�-��ӿ�~N�_�4�1u^7�wF/�>�v𵀀�ש�3eKU�'8&����y�uA^��I����V�"�U�qT��)�=��G���/� �ui0<���Cr�i��p� �SڌX����&ѹ7�X$��?���qza4�z���3�A%9d���:�*9�?f1Nz^y������^P�#�����A��D���9�rt�\hjiu��MQ�m�������Cc"�@��ܪ��:�n����+��,>/�ݛ��t��)���W| #h�˞��T�g�Y�J���'��#x��C��`��k�}�k�L~�X�f���t��eC篪������Z������	���cp����؀T��u����ק�!��r��_�Dg��?_���5j�yئG'I3I�O�\�ۓ�w����~��e�gI>��-1�b:ݱ E��Pu�p��o�W�w�Bߗ%�d��Jl��Vm�A]_�1#1X��օ%	�UY݇�˼�= ^.q̗��Y`�_4yY
j&�a�M�y߿;r��Öչhcjc
*:�/4be����q�/����c���am����{�ϊ�mZ�Ӫa��]�}ʅ���UI9�&U���`[��*Ͳ,˙�'��3������Jb\�T�I$���}m<��a�)����퍴k*N�xx=�������-�	ߝ+�0Y.�
-mV]���]qq1��8Ƕ�,&�4��25v�xZ|9i	��(�p5i�ѸZ� nK��y��#E��)�c��t�=�Kw��E���N�蹿d��&ۢ|��1�<Ey�J�K�˟��ZQ�[��M��&>�yٖC Up��s����&�:my��۩�|��A���V=n� 	Bu�����D�J>F��i�������{�B������f/u�F���re��`�?{��]�k�l
��v����
�1��,]���(��j 9�K9�ұz9���W��ᮐe�y.����?h	�*رM��c�"A�M	���F�V�!��)/�_�?��_c�ر������/����մ�CP�Y��E�
'�F�7tܖ��yYW괕 _k�,���|7=Q���g}�HCd���<"6�j�֎-�h��@�GBi܃��@����ܿG�$�
�4�P�7�A�Iah���d*��d��Mx>B�I�83��]j,V�2�X�^闊���۽p� ���!y�V_W��ۛ��˶ ��U�O�(�g�H�3"B�V7�1��s�\	�����c�s�?,��� �ps��um���.KbF`�I��X�t\8��H�A�ڒ��T���,���!�7D��L@�'���3��|3�_3��C�27� ދ�IZ����j�{�¬�z�q�H\����C̱��H�᩿��Pm{9��yd�����~�SP��qþ�4��6~�����L�Ւ��,�v���G�U�[%��y��p.~�S�j��[��V���'���׽�}�ʺ�������:|Վ���;�s��$�=o�"�z���
���� v�pG��(���]���:�)���<��Xp��;n?�J���u�:�N��6#T�0��2���]�ׁ�ѕ�/l�d̈  ���w8f��:1��9!�/���J@���:�m���Mqr!mBOofk���H�\zK��WT[�I�gM��;���v/vտ�ϡd$y}���)���J���72�SΤ�%u��4��@��v��@���Y)<�Xժ���^��fc��*�r�7T-��I���_}l^��	>��p=3�z����؁&ӠYsn�m*m�L�E��V5tēw� ^�]�$Y\A$��mL�=��/����p�&�q���)�P�n��ZlS�T�GD�Yc^3�1�71���<jA�T����ArP||��jFP�\}����R\��}��M}EF�A%�ʋ�oE�{�I࿹(-%=e[2�����ezr�����$�I�y_-�.#���2,6s^IZ�Kq��9d�(�K��~��m�5/8���@t�r��Q4��q=�da�E���Q/'����YZz_+�h\���)�}j�s�����tߘb�7G;���0'�o�����d'T�G�U�;�^CU�����r�%�tp����z6�w9��q6p�T����'������%E\H���
�g����Ҫ`�r"�T�u���#Q�d,��{}���$c�9 �!���+v ��(��6)��^��0N���6s�F7l�`s�ș�«�3wm�9��P���S��?Q�9�	Z\i�1y������K퉔@�]RY��ɏ����l�����6����(�ũ�R+zj��K���ƌ��63�6�*6t'D7m�G,.��p;
�S��n���׍T�.���6 ���S��A����q��}�����Y/�E�0����5f^0L.z���õ����Ʉ�t6̙�q��Ai�6OBiZ�į���?�٣R)5/b{������R#bH{��[���}�g�E�)���V�!bq6�!6�v��!���#�m�
���fTN�r�ߖ\��<ݰ僽D��SP$Vy��?��+����N�sa�9���.K��
��Wa�ųV�V�p���le���z�8����#'�Q9�oD��ׂ۾�*����Qzc��a��=��Һ3t��v�娶�f�^\-��ϧ��i~4��!�gq�v�0�Ճ2�b� �#�L���/�8g4�=�����	��W�|�~��7.-����>&B��6�ON$��T����Q"DM�Q��J�aP7f%��@zb���nM4ɓ��}��;��l�t����z���l����ݯ�͸
�@��R�t���C����O�1����	��g�{E` Qһ:���`�]��P.W��ڨ��y=8��̭ɐP�n���2��M�_0/�
�=��W��^TJ$�:��{zE�U�i��c��J��ю�G���M:+Fy����夑1�y�x�}���3��O�Mt]�>xߑy�
�B��&k)Φ��&M�d��,���3�6e����9�&nW�a,�H�0g/gy���[)�HTy�J|	��+�:&�2?�*�7	U�}![Dt���l���Y���>߬�E�%�%����b1L������YLm`�c����T�9�"OC6t���:�F�Ѿ3�D<�lо�~��3
��,�ՍU{]��xi�l����T�� ���n���]b!�$�i VO��3+��Q�*�m#W|���x����"�TSE�J�V|~mJXJ}j<�	HٻS]1���J`�W]J[�x�q��mh�,3C��`�ԝ!�����:��=|���/Э�E��;1T>���������V3 ��^�e���|�C<JӂD�*�=�E����'�u��rM���*���<ut�y9ˡF�(~� �v�����ٗ9P��� ��d:���l���W��'bYݛr~��_2Ԕ&��6���%�����tmi>놳䷿}Q"aO[�w5���r:
�
�u�@��rq��U%(~[��.,�%*��o��L�
���\�w�\�a!��GV��%��O����|fУˣ*�^
�`ؑ��"��Y���ʵg�3&�X}�]�֯utFQ���*&��{U*�w��U�5]�̿q���|�TN��ZO�E��4��Z����4k-��Di�����n��AI�ʻɒ��9_� 卧8.���#�IN���ؕ�{�S��5ޘ�OcSX} V���%/m�dZj��V�d_��M���̻�f��l�E�Ǘn�nP�Α�*)���4��.: ��]4K:����ko��w��)*@����cV��z�pD�:ت�aj�]7� :l���o��yY3����S�'����©�~�v�Ty�a�:bm>v�	���������k<M���CXf����*}	�^=�[�`�V>���&�ߗx�ud��ϔƏ�~�P��<���HC,�&��Vl?��tS4�Z�Io�,����M�b���!�s8-��]�fe�<��Kd+��Y�	����
�1!�5oSl�����8���Գ���K˼KI�y�N���E���x3\���C�f/���nLx�[�����v��.�xb=V8��7{q�:�N�d�����:2u3ty�kAOƱD�E659���0J�e��H��<f�[��-}�	�7�[*KMg�8%�)�!���v����ߡ��R�����q�Zdvw��
����E���=�o$��5U#޼�u�3|-��~33����wc����ݷ��f��I<`j_3���T"���B����mk��b���5�Lt8	4�E�%�ヴ��+����b���e�*x��G�����<���C�DL�Kǝ�a�T[sht}�$?:6��T�-+������F�z���0Ӂ�A�ȩ#ޭ��4�Ar)��AJ���3g��`��o]����ݷZRo��f��i��b�a�	��I��r[��#����%��,��[�m�߯]�9B��b�f��]|Q�"��=��D��t�E<��->[N�m;��B�U�������Ug����r�c"@/-�i�=(R[�"g�rBG���$��=#y�AOUK�;�8ן%#��718�K��D�,�F�����:���b��_���u{x�G���Tn�1򌮎v���Z���Z�aѥ��ٕ;�Db]Bx���γu�O>[(F�"�mM���`�מ1K�s������ٔ��Z����7���<7�np�SN�s���W�D���3�eK
<K�_���������(�]�^~�+=!OP ]��oh<>}�{�$m��k�z�4�w`�ԗl/�1�"�$���%��ه�w��+�{�;���'_��BBzJ����t<��e ��A�[{q��c��M�/O�d�ע�фw��hX������6%Yx�K��S�x�ڈ@��,b�oY�nQ�I�Fhh�؉bE�3����]/fQ0��^D&f��lhV;�����5��y!�wI@�a�U}�)��i@����E��KY�vd��X,{{t�W94a1���?\���<Y�e|v̵K�8�������tc��&�%����h:���C���;p ԰��q
I]nV�?��jz�N8{P�wKV�&�!�M�<:5�.�IGk֩t�p�XnIO�c����х�wC�tO6���֮�#�fqrJ/��[�a�~Qۂ�l�qV��}�wr�� 3kz���U�ʖNO��^�(�����+SLD�Lo���|�D���gc\�d?ftS�R���A�Ě�9�)���U�z'9����լ�9��N˲}UЙ"���yR!�қ"e#��K~�[��ָ��#'F���<�SV����#AE�% %�U��	�~Q}�d��%Tp��S��;S[�a>��UȠT����+��S.I�}��D�&D +��]2\6K�<�jRz�k��
�Vm��)�%����\�����*3Ʃ��S��2�� �C�P�I�zD�Z���ZUf�@�s���@�O�G3����ێ�~����2��}�jB?�g���B�V���P]���x]�@8UnE�����z��"�۟�^6z�CC��)|��"��X�>�3�$��R��e�6t"���V ��{��{z� %	�UhkYI���ɲ��+�f���J�/Z������|��ɇ�{ F JNV��o+�����e��H| ��ݢMMWe�E7;(��+�G��{p�C�u�j�O�`W�ك�E�e���q�s� X� 1D��T�T���1G�� �œ�~V0��cǹ�S����DJk/]1õu��4�QH~	v�@8,XP�It����k.̕yE;���}���n��Pe��[E����.m0<�NǙ����ㄆ���>��K�Z�u��\��d�*-���QV�D���;���C{򺌖�� �F�_�Ej�Z�#mT��J�p-�y9}~�+��9�8c~�{��'���0����0�^�KkV�>;��Ց�
�g�M�����,�@���� ԃ��
��ܣD�(���
�(��P&��-�#˚�7�,��J�5�j'�![H��O��b�N�����B2��*�3ؚ�o�IG�f�%ɖ�F�A�^��u��rqB�#]Z�ӿ���fU����s3D������]r2�����d���\m|SKt��#"��+���zE���t�ZҼ�E�.�@lġ�o��tQ퓼,�7{���Z��2��~@WY�@�ȶ7��p*���( �C����6A +lp2B����*e��p��T�}o�*������c�6g�{?�<0�� l0H�~�Y��"K?��[zgz�=bX܆߅��>���|�^�n�o�(*�����fM������Q^���z������=?��~@�䂡�u�";�SuP״���|x+Ҋ�&E��8��k�oy��$Z��սް'���6�>(e���������z���P���g��j�`Mo��М�����tԖ��譐HDU�P�n��kO�c��K��Μ�lk��Ew8��7>�p���=�I5�	V<1�����\!�Qpń��b�ɨ��OJA��I�6�!V9a)w��&��g�ޭj>�tYI,)�u
z$,q�9��ʖ,��E����gm"��aHk�y+T���@^�_���q%����$���\�p��3���ȶ�ܼu���\�~���b[�W����[��9f/���TuAE,��Jʜ{t���Ѫ�Uh���t�w_�<{9���Ek���g��5?�2äq{ء�>1d������sDحh�̝��-7,n6��U�J���Y��Q��	;��9�m&Z�;������]��l����i	u�SA�3������ ��׏?Fد�K���A�s�B6�f5���6 ��C7��	��/���'A�����eo}s�cu�[��G���.)r<FP8)��Ȼ�;;���-��m��fH�[[��sܸk�5`Ern���"P����]f4���>u��A�����M2=�������5��7_��9��!1�(O"j��2ө�-D�?7�-�m���=�	�W�>ͩ��|�]@�u�,o�bObXL��8h�LR��4kyk�p�^N7�$G���Wo8�=�����>Q�֏��L) T���2+��t�d{%��x��9Y���hj��v9��V�d��2�X֎]g�T|a��]�4(t��L"��|���c�d{K�8=<
\�ߖ��-��ڟ� �X�khUg��i��ރ�c�QQ�.=B�'�:�R�`)���k���'� ��a�Ë;��qk/�h/R�%�Z}����"�]$�A�p����c��L=��u3{��'���d<�7@�� �D ����Of1���C��?A�|�rz�f���#�{�_1���g=2������x����w���9���w)Ma��ѹ�[������m4��rnܸ��\M�u�.�T+���]�D�ј�	֙����-@6jYy���l6 ��L�@{�������&N�3x�8IM&^��j��4�(i��'�Z���D;�h"��I�H�4O����������RJ��W�\4I݊�wf��W9��EeH��+_��jRw�Z���7F��,�N�hX9[��)�C��8n\������=0�n�]�s�$�;
�%��oWB��e��׽�Uf�<��5�aIL�Y�e�k,�i�L�b~rf͖��&���'D+yX��c�U���o[���y,[�Sl3��7�wҁ�W�jn�I{Շ�b�ȇ��&ܶ��F	q˛V�Ô�_��z���ю�7���=��g�q�� �籒Y������ ��9�Im���? ��������HT��L��w:_��O��<�kpx��A�ێ=��k[��>�o����ri)��$t(�<}y��;0���{O��%��`*7c���1�WM�Z�����������݃C,��p�x��фZ�	�6�-)v��K:a	�݈�o��D���g�'����h)��	����0�����B	j$��+���]�x�N��u�j��`:>YK�~�F���P���� ��4��]!�lä�46)����� /�'��\p��g7O�����$�>j��y��:Z��<��+�5I�W�@�C�M�7XB����B�eO���W�!u5m�JZ�J�/5��M���V`f���y�Q�x}���]��H�7;�r����*w'T�U�-x-�P�?x��t��x��BV7��=�i��b��]eN��@FD�����ͨ)f��oL��<�2�·=^ f�����Fo�&G��%9$�4����r���k���2vd���c��d�V�֪D�x�󲋆�^]�#�tY���}X�y�bWa�[�0!�#M��d�'b��K�� ^�����Wv�l�=H�C� ��[j,I���u��i�.Q}�-Au�զ
��=���1��D�Ө*�Z_��_$ف`�P�n����3��I-�R�����Vp���8�5�Is���F�ٔ�1��W�Ș+{gs�V�0.d����M�ӳ,<8b]�Ǚ��8��_�|=e�)HT��T�
m�����H��!M��;+	W�%���:7���&!C����%��˓�^�O������5���喨|�%��C�%�݂��� �� |��
d^?��j" ��������s��ت}4d:��o�)���{����r�<TS��F��?ȫcq���+7��te��W�������B�e���"L���0G�OmM�=@h�/Uh,�ۍB?�ҮC{��ZA��1��Lܮx��p�3��hr|c��Ō����q�j�E'�^�o�1�u����R�[`i�Nป��5����R�R)���6M:���x}���������J�̉��3� �gA�o��w���Q��u��v���(�]���Y6��Y���WI�p�a�ZG��ڌ7�Z�^�h�7P����)��k~i�ڇ$��L������P�e;�&�}�'��!�'>�c>j�4m#�(�`5��/�<q=,�\�qg�]m5��8׷����+�>���	�|���OH! "tO%�Kƨ7YT��C�W&�#b�Gu��\��^2M�_F8��RRMz8.e��#�
e	�Ik47�wr��C|HW>�ާ��>|�m���h�j��L�}��F���7Q��^e`*�'+�0J��q!C��\��XY�T]�3mK�0T$��S��5U� �2�p����~���d������}��)�ݪa��w�&ч^��2N�#�NМ�u�Q,�M��i�C�/�4N�{±�V%I��Ӫk{X[6�u���q=��@��]4��DK��d��)��@3��D�La|��J�\�_	z-y�2�����GXN�r=��qhI�g�m�����!�rğ�N*�����ڦQ5���@�{���oӞ�i�PB>�I��(r9-��nl�=\�r�P>+��?$-��;�[�����qj���]�_*ۯ]Z�-�"T���8x	` �s*O��y�C����3��B��ӘU�[�/ͨ*Fd!�Ys����M�8c1p�Ȕ���
��$K=]	�}ı���A�u�H/����<���CS��E�<ȣ��簹�����'sڦ[��L�#�w$�����O�P�ޯ���nU�P?�
��e��t*�������B��R�*ڻ1e\ͧL���Xɖ�G���I�-N�T���%Q�<�os0l���Q��sMv3���c[�K���J��U� rf��F��'Ջ����N�/�ԁ��i$f@Ӻ�Mz���C�%��Z@�?`����1쌠�+IQqM���a�.�FS>�/����u�(�#�K9,�W�!r{S&��a}��E~�����+G� �{��f2�[�-=J@+��F�/�Hihi".n����W�2���迻�X�ڲ2���cѹ�u�����#�5�KƀF����#�a�*����|�W{(���4"~���Yر��"�?e`�l<��J:6E@<�p��Ϊ�7.��'|�
�st+�u�螛�t��qT�c��&B�~;慝hO�؋&����ƣO
�Ϯe��:�r��?}�-*W��T@Y�G|��]�t�}y�e��?�B5��ⰹ's-�fة�D'v�>s�z�'�K���V%��k����D�����)x7�c�.����E����Y����˶ǡ�nL��������٨���=�K.�cQ[�u�jZO�lim��A�M#�r�&&C��E�F4.��,�ظ����]h
�$i��(��I��;�`�Hr��d�)�t�l5%ś��@ak*��n�+t�u�'UAI����b5��E����IH���A^:���A�>�~N��G�bNU��"�.�	 z R����)P�,d"�Ԫ�b�X�e��U��$����3�����P&��ii&a���d��s�w�����X����X�E�$$��.	�E8X��2���lD�]�O�ޜʧKK3���2�4B�ω��U5n(?��@�W9W��Ie��@<���
�T��ښ����)^e>i�4)�'H����(\��������"��_�@���;4�9_��c�#�V�d�s�X�3L�r7`)]��6���s�?ne�ƑP����4-��3��o nG(OӌMz�u�����蓰6�4!Sy�S��c�����Q��s�f��fN����@1v&d�~�TMry��ŭ_��C�L�Xި��!w��79]��K�Pt��Ft]���h��R�*$˿V���{�a�%��D,V�KlN(�8['K�5D�6��-Ǔ�%�
�SYK�`���׼�U��#�o�6c����M��>'�A�1o&�{��2kM`|�0T1�9�CN��t��(,W�)S�]i�%?	\^+n����?	�u�֬�a{�� 힟����:F}�y:����>��f��(?��8�o�k4�(�s��ٵ�풧0��Jsұ���v�n(��z���ȶ����6[����Hdԕ�j�g�n�C,�� ະ�%<>���P��c�"��Nyǆ�� ��bшc�#���l�{��%��%U�}���QyZ7��2�Ј��k&	%�ty�[��&�3-�1��.�\46��)��ڂѐMe��x ij�:孍�-ϰi^��*nl�8daaH]	����Ldh�r��I���2�6�:���8��0v�u�E��"�e���b�۔��,8gR�m&�J:s����o�dSY,oc|6���?��� ����x aNC3Ix�*2����B����SQ�����X:��D��\��1l�i�y�v�Cߠ��������#+��=����n�~I�5��q�!W�
������&�S��`�h�&�`FI�\��OX4+�Ѩ�-���jѼ$�l��Z_�}<�#sS�Gq�u����U�����0���d�+1<|�cg
@���/fL��[0_!ڈ�u���d�d<[2çUTNu*fJC��kb���9QGX�� ����U;3;n�ar�f@5��ʺ�7�+��A_u���7�q��tr7|��MZ��'����8�!$���k�dF�B�Ɏ>���Q`��( PS���:�Ou�T�Zk�c���� ���-�s�� N-�M�fQ�1i:���̶S� &���^���b8�5:f���jp�m:��7~�9fd 䩶�J�s�)e�i�J���|��M��ؔ*ɜ���K���Ln�Qg���y)�Xk5T�;���&���~�!Śs
	�1��6	sl[<~�4c��V��C �sS�D�>!"Ӕ7��Ө���0�&ܢw�I�����QN_�)�ЇO�/�\߭9gq؅pZ��h�f�謔��]�}b=Bk��!d��h���N��pu1��
!����ifV,;����G����ۘ�������3@����(BEN{	�����%��%��&lG��K��9�=/�Njy�lĀ�|s��Z�]��V#k�>��@¤9��o���	7 +�����}���9�T�`|�l�,�v�ݞ��q�j#�,�z �CVFt��Y,6+�ʊ-�$\~�t)1�������t����VQ?|�~�#�O�b�j�?i�H��|�h�MK��M�X��B�A�kB���t���<����N�~b�c�P�2x�k�ci~�Fck�aH���b��̪�����-j�B3D3c�����i��V�#Wq)dt�$\��*)O$o�r(
&�[$v����I
�hTY#����<L�i����F3݃�z%��<�l3�8��}.|�Y��M��H6Y���PR{O��;���?�����66ë �/*:T��]N��c	'�Ul��z�� |�w����
�CVF���� ����\H|�-T��$)*'�~45����!mg��#R��nI�������5�Wy>�cra�/)ȕ"A��}M���s ZF}���#�������� ����G(,^s�|�Ҷ�����=�_�H��@�(�t:"������s��4�/b���9`��B��a��W�YB{?ˤF�����D���F��Ƅ��	w,?bd���C6I�u�R<��_.*yE�.0��FVi�m$��S��<�q��T�]�)���q�/����P��=7ֳ5r+4��]���s���j��>������#7`��֑�a�J���F�~fv�7�k��[d���V�Y���s���^�&������X��s6vLA]����ψ]쇡O ��B�߳�πZPGҋ�Z|k��	�)�)��C2Bs+��ו����a�����>f��똬	����{k\��7NHÜ�H���2��B�VC?��K`.�}M�Ϟ�ĵ���"Ee�)�Qߜ�^Bp��,3�Xq}p���3��[��"�9�_�������]��L��׍BC��?�ݷu�$�
�K&,�eyS�f��@��7��}�.����M��]|uԄ�l�<@�j�Gz��W�����-���D�en#�1�mbW�H�Q��k�c����f]-�ѳV�ˡ��EkY��z�l����!E'�ln���rb֖�m}�������6�2�D�$+͏���T�3��a�V)TT�h'l#��E(XEt�[�T�,�V���
A�ҘT��{ /���ﻳ���t�6( �7/�`�� �>�վ��ױg������\˫`�V��6�;h�,YY�rz�x������湊q��� �n���X�x�M�1w���7w���.�u�&n1C�|/	��Aظ����"+�l�$��EN�Ϭ�`��\����rs=n��+
�S��b��];��j�/k�8�a祝�K���i8E��1��z�A4��%Z�����X���>���ᑛ��[g�(7a�Y
�0�*{�
��,����SHXD��ӥ��9������������'��\�*�{[��n�mg�x���� ��+`Ӣ�>L�H	������\�V�q&��S�6f��%҈\��{�i�@���0�k6]���S�8���yL6�{��Qy��D�ء<uh�G�e܄H0�U���(tE �c���?1<�3��`�U��\by���D�X��q �]�D��'g5��T0y��h/Qc~�	ӑ����֟���8��Jޥ����?rvLf(x���'�+̝;O���$B��	BT��Pއ�	էu@ާ��u�����u���A�L�i��Γ�6�	s�`�q�^5>�.TUa�Cly	)�-5�b��ޜ�S3 Q߬�p���z�#���[\�1� ��Ut�(��Xi�}_��o]T�!)�IF�?�͕�l���"fz���4��|����,y�.�f��F�j�]����gΐiL���T���-?X⠩�|����Y��W��$����Բ�~_N�-t=��c�>�5��Аi��P~-�C��N�z�Rx�}Z��EfA�2�5��f���;��#P����*Y��k�uR���H�Izi���@��ʯ%]���1j� u�~e<#�����7,��!�@8�΍�
�@,�1��*�rS�!�rJIV�2�5q@6��qi�f
���������6O��*�]����)����n���8��n����ʹ��uj6,���q�$���!�%����.����t(�dg�x@�wNO*��RQ�?�"`��`�/��@��ˢ 4���b�H����1�t.�>�lЁ��4�$�Z�k+�IH�x��1|X�= }3���N����1�!����d�xƖ��Atg�'��N�O��G����?�>r9��1��6�L�)ǀ����u0������bke�ࢴ�a�[P�Ѣad���E����	'�IT[F�}G��b��O ����
�r��P+���iEG	#�K�c(�@�b� y�����	��� #�sH��\��?�HR��y8Z�SnJzqif5v:�+CgS��f�U�_��Y'9���/��
�tT�]Iq/,�{����i�l�!ͩ$�͕�9�d�m�;�~ !�]M�pj�N��\|&Y�_s�8�����_Q�]"G���͐ޙ�A���d$@�2��]ny���˙��u�X��d�,��Ql�(��t�JT��=�d��7tj�k�S�	�M�h��i�g�������	|��۪�R&���Yx���2�.^j�
?/N:���xmO+�=�Y�[���,Zko��r��K�������hڌ�z�i|'^4�j��
n$�T�>�%f#����9���	���@'�Q��d�_-�&diC.A$�즪���>Xt���~�R�o�w�3�j��FL�V��ED�ȪɊVu3�q�2˿Tb�(��:祪��)�V�(��mo����9cIR�K��A��_&��Q��̑[��I"߳|H��^��_�R;��|Q2�����8|�S�{�ex��������������"$۵ˌy�'q�_�ro�Գ[U
��"h���#�5h�6��zZ�)6��+�C	���ﯮ����o#��<଺G|�����3��Bds� $u�	���8�a��P��gUm��~��۵V|��}��������sLaf��`Ǔ~�u3��y�H��ڔL��|�����/�N��S\e$f��]D�F�S���+r-�u	���+��L�����7܇�^kT���R:S�>�eÏ��RN	s������ъƦ�w�̭fJL<���-h�]�ڸ��ދ�緄���#�r�&TX��UgD�Cϛò�CX�)=ڊ��ɭ����g�AJ:[=Osp�z�^�	�GAݦX6�7Ho"�D'��v�3���0z^�:([ꂩ -f�H�ma�K��&���+�]˳.	}XD����`��+�y~�] ��6�K�sܝ���:c�:�?����-.@��� �8P�5lp�ϼ��PN	E���� R&��C���CQc�c�'�߁�:��bE�v�8�ئW��,� �o	H��)>f(w���p[e|�`���"�1ZF�,	��e�g=DԽ�@��>t�yV��r79\�s��FQ��U���p�×#�!hQ���<�%e�*[ME�*�pxn��a=�Ӑc���q�w�#!6u����#4Bu_e���׻�����P����{o�/L����U���V�\�4i)|�4��a;B���>��4i{���}��)����N�t
�z�q�q'�K�y�`i�S����ZK�Qj(F5l��>��=Ä k��[ hS��&���Z82��c:D"����q~�BB��M�ZbY���:נ�#g�3��E9_
�5)�b��Zc��,�L������� �*��P�_�����9�LpBh�\\HҬ'�`��[�b	����w���\���H(�#iอ�Xޝ�Ё�0W����ʒL���)��/m'gW��B�(B@{�{�bp�@)f}�W�����^���I8e�U�sh��ǜ6Y�zd2�@�!��mA��M9r�AgQk?d
¡����.�X�&�(R��ɩʭh{�B �U�1q�/�d��<�W�c�(�D�[�V�ѐ<Ѕ�d�eϱ��L���u�2{��y_@�jkS��OJ2i����QD{Z	_��^�n�~�щck�4 cL˸d�|��p�Tݻ�w�W4D�T��,�O�ҺZ�K��O���K��b���[c�M��W��*ݢ�1q����ay
b�B�	�Nf�ќ��GOGKV�����.pҳ:Q%%�	KUPʏ���[�����(�j�z"��@U�����a\�mnl.%z��0�|\�� ln���`M�MᢚǟH�pI�Ї��� 
Y&���Z�����o�Iʄ0l{��"�q��oT�7�tfg������p1)�ݝ���q��kљ�g�/��9�)Ǹ5��#ӏ�|`���������Qa��kW�/\�3�ĝ_xFM�a�W��B�����_��9��j�5���'\��Q8C9劚�E���6x"�$q�_�]%�y�`���F�ex��|�,�)2/�K�����I�9=���D���k���!PӲ�R�v�dx�'H&+���(6L���s߼�怌T��<��@��L�W5�� l���W��>�6J��i��[!m��w9\/w���KD3�=ڍbd��FQA�4\�v]�����}W'�zr�����5���	��3���lI���&���?$��])�1�e���Pȷհ�ֿ��>��B�܌�1�±���9��ErE�K�N��l��2�C�r��.��^�ɽ���b/����y�?�D�z9 J��ƥ;>��&6��4�'�,��T��̚H��(�"��f�c�*%BXM'y���QS�J�g'9`�Hy�w�ͼ����ɕj��g�M?rS/������ri��,�$|���kZ���x�Ӷ��"ԣ�<�ת!�qįeǙ�
�d�cÞ��B��e��!J���A��yϔN���$݋���{��oxvQ�D9�z�PD��&h�Ag�(lS����iX��N��Y�jU9�I�W�f�.�Gl�-��V�[��FQ�6�m���y�����������Fz�j[��#ҽ,��Lħ�W}��_>�������ȓ���招�� ��}��~��2�Bޣ��o�U�l1o]���a��L���5h�)�5e��Gl�P!6�h#bH��j^n�_�<���v�*�3Td'_���6�d�	[�..�2a3�ϛ]�zF�ο4 �v��$&貀�,L��C>�K,� \�CG�4wsM�0}���h�~#	2ʯdԥH�I��.���TS�F}W�BL� 'j5=(����%�=���~3##�f萸ݗ��^�Z�-��gCN�8��,ӹ�p�V�}_"��<EN2�1n��3�h����DvР��=/a�w������K�E��]�}b��)����X	l'���x�n�Ҭb���(r3�y�>��G'9^�t*��MvH*ԙ���R������]��۞Y��vq�Y �SP:9,9%gľ�����ʄ�+�"�26���׹.�+�M��U�I�"Ͻ����R���8ށؚ��_���)�����vF�{��eo7���)L�e�Xҷ�.t�r`��R�+)�l*�^�u����`��¯;����!��}�Gd��)c�E�4Ȥ�0U1�i��B%�׀6"I�'.6���H�y�f�s"��{���r��>�\��B�u]@BLU��@�b-�:�Ф�C�)Xm�����ioR/��g�8�k�|MnT���l���O>-eo���ϥC�W���vö���_��d��f3LqV�V;�|C�b�� ��=��У]���L�r���A�ƥʃ�f�M�&.�e:�_�7V+ӷ���r�2�E���m��l�¤��#�ŌgS��(��%��*ي�gޘAgiM�6��%�����.��O�@m��gHp��69���ow͹��N�w$��?2�pF�	���H+����`@bМ�|>�͇�t�SQn�>�̙	O{ɻL17�O��T{�����dW�ʹ���L�/��+l�P�'��Q�gF9(	8��p�g1�U��Vpf�]��
���#'��G�?k3R�H<@̽@ue��)�Ȥ��|
�����T�r�l �����[�]l���0P��K��#��$%���?���"t�s�3i�'Kں������9�?���'��`�	Б,NR�����S�e� �8�Ln!c��!�ǯ)�Л^�)7ԡ^^�d�~6������%�������ߋ�Q%9�1"3h���d#������m�p�2(uۖ膩~ʙ��MtE��@.m)�K���A�z�\����{���Ȫ�|[����$���n�^æ�-	 /̋��d���ʬ���u���ax���ڪP+���G�Vĥ
�^���i�n����A��N|��[���c���@��C��+��m�j��Ee�ܴ��S�$w�J��Lv&�}���uP9��u]R�^t_4��J/+Pb����9��-�5���W�-WL�b|d��z�;��?���nE�������~Y���"H���򄾻�eq�$�2:R|��l�u��W"��q��t�Z.>w�:�|�ןA?�r��O�u���a���j}0ϝ�=��	WyE$څ��ah��C.�2\�Ш�M�Y�V��A4W]R�AuEh�B��� �p
�r��\Q�b�_�e���F8��P������p�Ũ�� 0/Jq��iG[�P&��(;9�J7d�G!K��8�p�Re�L#�|���E���:�� �K�=���Bb�G���oI���ƿH�h�u��F��E�olee�y@�Ꝑ#�fr1*��@>^pwE���Ct� ;�^�$�!h8f�����)���c�X!�~���g���w"؃:��G����b�E:���}�aE�C`R��#ve+�K�0��H�ږo��j��3�8r�A�M�}g�bs�;��W����3�+� �z� \��d�E���p�9|l=��A{��W�jc��ar���ɖ�i��ǿ��5A4ĺ�F
�W�N4�J�y����g�����Կ�=#���_\B�3�P^?�3S$����M�A����R��|�Z�#�./,3��V�B�nɳ�M^���q�����g��5��K��A�(������k[��dc���zJ����5rK'����ї�xkAd�P�C�L�nk�$wX�G���ש�|�9���|'ʩ�Gu�yտJ�]0��=`d��k�.D�,q�Vs	\�F^;-������Om�&fz�P�<G'�V�K:E��l]}�Q`�G�
�øO���a�jsBcxt�]�Vp�Nv.z����n75��D3��4}*W�7KK����X%����^-
no�=({f�}U:@si����H��{yi�62a�>ĳ��`����-Mkl�wU>�#r��+)E ��ЅE"�Z��W����,�[�i�Qv���+��\{�2�Kk����*�����D�g�]R2�q���B���~r���©`����z��CW�AJ���8}�'|�Xؖ�V�KB��M��
�#�Q���`(PIjL�*Ͳ�)���p���W����N�����[#=��A�w��)���1��6�އ[�z��R�76C���b��D-�i�ݒ���m_��*����B��Hk�E������S�9��?�>�ό��%��wZ�n7qn��-#.p�F	�f-)��{�7N����',�dO�	X,�7%�cXU��D�D~Le_$_Hxw#��r;�B����Fw�����9D_8�R�j68�����D~�����AO+��4d 5/�!M���q	Ӌ�߱b@�2��9��:���l����B��첶p�j�4���\\Cco��:m.4��KE��6��GXv��1��@3Ը�H~ �	��Щ��QOsu���um����0��� ��XR��n#�7R�1Q�;N먄���!�����y��Zu��uQھq�4�.��&��m혹����d��gV���=�DB��s���H�h���ԡ��o.Ӱ��֏$�c��^(��� ����4G$)�=�����vb�B�	����M	0e�xt9��QqlQ5K!���nv쪻{��+�3�t�����|�P�݆)�(��dQ���7%��k]Ȕ��0�7��5�9Qް��+�葛#��A��V\2�E)�����$�2�ʖ��X��:_"�B��h6�?��>k��;nD �j0h��=;	?���N�J��ܩ��P��<q��X�ߡM��=��Ri[v��"�<��5'α��3����ˍ4]����H�i�bl[��V�]��ꉤ�n3@���W/55w'2�l� ���,������ep.z=�(q T��(���� ?d,QqY=�Ϲ�Zh�q�\,��^c�yB���a��'���4��;�\���j���HCS=*l���.EdG0����=�P�~�nX�
�n���by�.�{>��&LȗT��f�����,�!x�xZ��FY���TϷ��A��h�ʩ����ђ���?��o�.#�����M���IA��J�!���*���1'�iT-�Ϯ;�Z��0CV�1p���q ��A:����)���XQo勬�z������{ì�C>Z�FsUf3ڳ`,xr	���ӷ��pjK����05Rg�d9�ESG�k÷���Y�}���3�ǆ������<��F�(G�rhO�"��&�4�☉-d'�S��"��	����bζ,T�e�w�����E��d%��R{էku�GL%�@����I��o]���kP(��.�[^�0tZ�Ija*��}�ٍ��M�ԯQ.�<,�>�^�c�0���J����ێ��\�
�+r4�,˶W����h�ѡ�;͝�ǵ�,uS�ؾH�^� s�~�,�:�j	rŉ���m���b��WҾ��/����)�(���/��u�:o������ە8;~{��E'N�!F=��� ���ݷf�ק�2|I�첽dϚ�|��i���?_g��S��м_�D��VXpn��,,$�{���S@ɏ���~�`��|�M1+Ufm�ȭ����)�HUE�k�������7�c� ��K�	��������a�p�Z���Ѱtg�Ie��E򛹇Lb6֖���沑dH��-�7�@�*�k%���^�P�7�9�b� ����w�
G����p��dm�Hᦜ�o��9-h萯>"�yd�Ų	�p{��PH\�Z��7Ï���d ݟŻ�9s����~Jww�?o]���)˃��mRiC����}��C���#�xX�j��e�ԕ=9����$�X�"D ���x��3\D��c*lo�R����
��N�����B�{�0]�4
�f�yJ��T�o���T�Տ��E�����E+�2wۗ%�I�G��^�T���T�q�P���QA�ܜ��;�`�C��>,]�o��2X[���RQ�u���R��e��Ȑ�S�O�좠f�K>�Ea6IS�s��W��v{9W�80E�b<BLE�m�C��Et��<ו�z����c<�����B��t���U��
�F��2wm㬃����;��F���D�~~��V*���^�	��'�� �@�ǌ@B�'T�Q�~:F���.[��|$8T$ ����Q�ޛ3��/��G�N� ��)g4W��)�K'Ŵ#+�L,�S��"�(��e��gF�D�&w��YB���Z�#��^����%�\�&�b���Q\�:Bތ	�}�bɂĲ�D� |�UY�Rs���GנA/<%v�e2�7Kyw8`�XB�\-�	�0��+�R^u�7���镃�e�	 �,0�z��G����|�F�hpd"�ln�S�Q���=���wܲ�l�)0=��׍�H�in��gPǩy� H��7���������B�1R�%N�������D�f�A�ݼ�K�ԙ�۵x�H
}X҄'u�0�V�j:r)5GT��u����y/���CA��;l�Z��M�^L4-�6u����� U�W�ip-�5��=t�l`�޴t�%ƣYqy0���>��uħhZ�8�5Jh�^�q2Q���*���8܄`Xf	��S	���wҰ>O���W�ʁB(��'ٕ�e�e�u�u�,l�#|�6y�y;|��3��5��&2S�q|�x>ӛJ��s7�0�I�)�i�o骗
v�Zh�"�w�͚	�O@�x���)�HcM�1�"d�qe�����E̾�;^������+;*P!���k�)mT3�x t��rpH���.�w(n�F�g�������H�w6���?�y��q�T��!�TA���� ݀�q���;�=R':�?K��D��Q*5�H���
Rn�L��^���`�ה�sk�������]��<�G�h�!������e����]
t��,М;��Ŗ#�X���v\кM�t*����5�hZ��"����q$\FX0����1Z\������{D��)�*�
`lBsǟ/���M�ҡz��O��xXj���L�-��¸�$������� c�,@3ޛ�Z�B�X1���==��
�m&gb&ۨ��1�|����e�z��h��)H��m�-�&(�)Q#,ߣ�=�N�*#}��=VЬ�fo�Oڊ[J{���߄՜MP�=�X��E��m��h��h@��GFr�K�ގ#f�����,���J198s0&� zU�.y�� ��E�K\b\�1o{��z\��>���T:���ь��_�FE������-��U��蝴.?�v�.��W��~���xIy���~9�6/[�+��&�Sj�0�`�Y����
���=�[����Nw�&XZ�ܡQ���MCH��T��|%e?���3�']�q�~����b��H��r�~�Y�_��k����:��"R�9��is�(�6��[s�y�����:�YE}z����m���#�aġB��z�~�����=�̬q%���'m
E�9�'7n�i���]�<��q7�.�Q�ʞŝ���ek��B�F��Z��/�O1@9(ȐS/���� S8�&,�.����5��+�U����q�v)�1�5AԸ�a�C�������w�����0,0�bZ����+ĶlWu�E�ڳw&P��ʕ���!��1t!��3p��m�&�;
��%�7�K���`���Y���
����
;@H�%��1�(c��7
���KX	EI��Q��kh���E�n`D�J���E�K9�}p.e	4�>�񀅨��;����3�)+�����>4����U���2U���^R�~�t�zU_̛R�|ͣW��Lw���tN��
��X>{%b;�3��erz��cB���1\&=�
�\&;b���e����g��:҉Ŭ��m���=� ��f�<�o;PG����['��0<�KS>���H� �u���f깺�����?[���`��r�ѡ�1�n#w�=�Z�UٴD�B�-K����U�����p���ƹ��l��7s�໰Y���E�*�c�S��k'�~�wua0�b�Q�c�f�%l������@��]�?��ݵerV�m�X�!�W�Tƫ��./@��z�����<�!��qhro��k��Á�+��:���u	d��1��{k�zT��5
g��h��ݢ��9ZȈ�t8'o�8N�+﬛DO��at��dN6p���p���f*�lg�~����c�����A����
�o��k��p�ڪ�n��8
��U�N���	U�zT	���^�6lX;눫f������ggi��f8����3:E� X��ig~��K���d�-{���+����m}@� �e3�Lnկ�C(�
�ځV	�7-�uX?Q4�*��19.?�n¢Q�l\'}b"'�|�,��������wd��K�w;�\ �\2.& o{E}��#��ϣ��u:|��y�	��7*��FmhM��P_�L�*��kmBX�i�Y?Z�r{��,�������0�yι�r���U�=æ��_�Yz$�4XL�]y�.&Wn��]e���7��N�������r�>�!����ɦJ��׎������u�[��Bk!49tv��<�]�G�HJ/�giC��S�<����k��e�?�ND��g+{e/ »�_��J��4���3y5�LJj5�����k΢���D,�;N~�)Y�:�zp�8k�����>�� �� �wa@�zX�Bel{TQuUpѓ� ��������mSuY��2M���C�yh|�w�	x��i SAgys�~@qY�����>֗/A���d�F�gN��+)�����"��B���u
p�=����C��P%��� ��M�Vj?��"%D1�6����7hU&M�~�͞��e�{9�)�
��3}��I	(r,򋓅<�*d/}?� p�o�l�zF�?]���Fdӹ$ �Ӎ��S�PSzS�dBE=!�j�Q�����Wq�0��̳�ʳ���E��Yz�Er�FE[.�Ҡ����VQ��i?��kN����8D�kj��[�f��,G�b��d,��%���s�s\�Cy���dk2"<�?�k<L��1�`�����68���'�y��s:[�oT�A�5��vkU;N�<�B��_�#EDx�ⶀ�
�� (kZ�0Q��h�p��Y>3�/�j���N�$3VSz��O6�r<]�9c�^btդ{����HX?���63��`@��^~����څ�It��/DY?��h�6m�/�S���3?��d��ͤl�(��ZP.ԈI�Ce�<�S�[�E�ZK��Z�MC��;�U����aT�nk~*���ɩ�^�ؖ�q���@罾��$O��K��ũ���D�z�xAd�,�A��ޗ�3]�������1X�͘Pҙ.���y�q$	6�vnU���&�l��d��d�5>��ƛ���＜`Ƒ��*�hފ�B� ��R�k+����H�f6fF�T�*���2��7~;�[��g��H�K�ʞ�����*����2��or=c;lܐ���J7�V@�{�e�YU��7�� M��o'�Io�Oj�S��HI�%�͋�yd��a�;-],D������9��C	)��@�Ώdr-ry���g�X��a�Z�q�:ރġ�|4�)�oy�m�^V�H�Q����h�ʪCЌ�����a�@1���Mۜ��ً����(�8���j��;�����v���X��r�����v���a�?~�X�6_XK�6=܂nC����P}��S��`�ov��[ٯ:��!H����"q�qG��b�pD�R�c%,��p�T�ǋ���!�ՙ�"�{�N�:H�\�iu����6C�������l�l����:W������s��Q�(UuV�̳�u:7g������C��~��j�$N�i��F����l:���@7-6����X���r�Ϡ��*<+Ь�B�0�ůY��-`�o����Bn���i�=� shV�m'�	��O���3����U��YC����~�����m}�+��C���{OZ4z�\�T�x~r=�q<�|II6*�Y:k�7�Z����##(`>�d;p+e�o����JR��w�?
���rg�5��9a}IE�#� ���ҫ[�6̝I��;��cK�Y�������7d��W����e&�;-��l�c����WO(7s�kׯT~��=����W�4��XX����;/�6fe� \ܣ��]ڴ&��;��	TC}��*��I+�z��ŤWGK���a��7�G�$�Q�g4��ť1S(!��l0��=��&ym�m��gʽD	�V���ߦ���/�
�&�D:N�?�w�{@�D�a�X})�=x�ӭU3�X	�DOw�T���-�ѭT���H%r�}�>�<���s��y^B���\PltTqH1>�V?�6��R�k�����b�y�VC�)�0���
 4jq�ǯ��彩���LQ���O�@�!4�Fw�U�.V\]~��ϳ�����(��t�H�.�p-�m�����'���`��t�L��>�>� �7�d���'��C��mQ!�h�WG�2&���9���M�N�p�xѸ�-�`;�W���3?���O}����u�,�u�d�я�pɎ^�E��YNHD�T�=���h�s�����[���QY�­��W�Q�sP���Z�F	��5�m�\J�w�=[���s�*���/K��m��A��IS0t6��n���8�����̘�C��/�6��&Z-�K*L�Y�\5�n"�_'R�f��T�ǱL��'������Ė��t�7�
�h�����M�M8�)�#z2B�@���ݟsiޏ4�Xu�3		ǖ�Z��ދ������ua��� Vd��}}( �ͮ͗�}ւH ���m�{�w�s\��4����3���ǣ��L�3�-��{ܙ2��0�$�L[���q{���xR4� $Cx�b���/{�*�Vp��"��ݴ�H�wo��h������d�z���2�%g�uo�0ܪ�)H���f�c����$�V��c�)
g����}�(h����/DN�!���nL�����G�a���G��lX!C�V4ns���B�Fu��h�θ�,��1�K7�!�*�q�ZߤǱN�{�c��wm�ڸjLeN\S��I0a^?�yU�2��j�+ ��e~��7���,�-d�G��d�0De�����e�փ4��ˉ�o�Z9���S`�>�׭�:���OK"��p2eO�]� ��6�V�;�B�I���o�`���=�֫흨������-:*��dl�4m���T�3�Էd/��o�w"�-�� #�6ߣ�Kn�]�D���Ux �W���Y
�3��դc�@�D��J����j�e�� ����e���5�����Ά����P������5�+��|��0I4 ;�"FM"���/�����<�a�����;�Kݰm=�ui�4ˇ�m�Б0�/�1�����ьCmK+�����:Wϸ�8IB��w&F�m�OR��Ro��[33 ��H.L�]\��S%x�lU�[�'��o������k�\I(�Y�M�ה��S��n���̛�U[�?���m�t�^�k��
��2�E[��Z�'р(h��z1$:1GюzDZ�i،m_������8�p ��Z6ԲH]��A�@>�X���k��1�of��ZT.qQRV_{d����;�ҞF��iX+�<���F�Pj�h�� {�\��M��G*���֓EZ ����xxOZ=�w̞j�<3�[%�Gȭr�<�Pٙؾh���0{�I#A�3S���Fx1��ȕi��Է��ح(�Ǟ�*���㑖5ؠ�
�H���?��/54��i}�r힝]��r�TM�*���L��[*���y$*��_Ř���jgxGj��d,��q�Wk��.�=E��o���aj2�B=]*P���՛����oN�ك�cfҵ�m���ƕN��K�m���-����]Ae��L�>�=-|�Tl\s ��|�F	�{���G��Ee|������E��㌫�@8�%�3H�셓��c -ȱT�Ne����<0���x�2�O�ۈ� %��x�0e�&Q��/K�q�z�{�[B3^���2�*Rb�E=�|!3#�M�����n�Q��3�P×��9��ʑ�
�֐-��Ն����Kǔ�^�x�@m����Q^����T~�eN�ceL%��J�O��c�Dbxo��0�eM[�^����P�[+�-�r��+�/[�. .���M�U��;�~,�-���������>�#�v�nY/ib��	F��Wύ�e!Ճv���o��S���x�ٍ8�� ���Q��o�SXhIT���	�&[��r�����at�Ci�̸�簊;պ��*���8;,���S�Ā�r�����L��1n��"�ȯր�4������Ly&Z\���:_U�56K�/���V�R�>%�ۻ<�O=U���EJ�r�pj���m�k�S����$���h(%S��`�=:&D.A;������o���@�Qf099�)����]��>;�3��Q��:�]���cF�# ��(K�Ժm)�(�X^H|��?â��i�Zs��oG��E�v\q�C+hPlAX��B�"'��T��-��l��J�E0�Y�c����˩��S��baLQ���TO��E����)��d�W"A �o���
�%�&M��X�6�fPԜp��@�w��_C�sl�Od҂�G�g��JF���xi"r�m+�F�v�d��2P:Ś\��Z���o#�';�Gi��[�`1���a)�I�n̥&oQ�Ya���B�N�ԔG��iz8��(wYp���&ϑ�����A���p14�?!�@�<Yo���Y�L����t!u�n�f��`r��͋篜>DgyG��H�+j�H8A�gߢap��[g�i�M��G1f�"�����ʸ�,�0xƝ<�Yl�,�#&N����	N��w�!� ���4�����C%އ;/�@vQZIĶ +@��]c�t,�d����G��V-Ug���]=�',�s&�n�Q'�n.������L��CC��q $�;�D��� �}0�QC���6�B'$�S`�m�4�OJj��3�:��c�e�¨�0{+9m�x	�p�d4H*��O�\�����f��o�}�����Os�K��VWYX
�
R&ׇ���n��#昱2���l�e�zq'�!O*�ߎ0S+�)f쌒����xdT���G��$1��ۥi��]�h^΍PI��G�Ԍw&J�����A�D���]�N�@���g��w���o#"��{Uv��^���7�~gO���C���%$&t)�9���q߇�T�>��#rߨ��8O�),X�r��@�~�+U��:j!�0�?��!|����٬�a���º��Mh�����������"IB��M�I�_��:�2��^ƙ����ETl�k���&������?�j��d�`}	�TL^-s�v� $�#��^�G2�[�	P��#jJ����U� �DH�Dhz�n���������z�㉸�kz�MO�a���x�l����!�wZ{��wޖ���bvD��yX����?tx�Ғ����'�n��G�(]�����{]X���'y�Ƅ��`��b������������;�5 ����fa�hf�R���Z��0�(�S+���M,�"� ���y8�[dC)F���8߶�������4Y^O��w�4=2d�WB�yC�w���QUgu�6L���G�
��B�A�9�L�>8����{�
`�j�n�PX:Ȍ���
C(?���p8p;�jZ�'�koգH���)��0�*H�7L�����mfQt(�b`328�U�3 �!����V�y�qu<P͗A�M�	�z�#n\�"� ̌5PLA%u�7[8�j�^�������x9�
l}R�E�՛]�"����2-^�kD�2���Hk� N�-�\񞥪���L	�L������� )����ͱ�+
K�]��V� �}"pY�O�U�� Qh{p�:|*�E�\�N4������lZzH5����!5J�m��.�.Hc����$�,�L�����'qB7�kj}o��+ԒJ
��nג�w��*��K����Z 6*��E�b�d�<�}�a��ݻ�_�!���+S�zվ|�[~t��DZ�����n��������
�/y�������Ω�%�8&�TCI7s*S�]��Kd��­�.�$/>��]�ͭ����Z�������x�}ҌVgV�dBm�{���*�e����!��Ҳ\�^ʛ5��H�>Z�+8���M�8�f�*�.S^0}�x��@p���m�U��S����KF�Ґ�j��o����Ѯ�<{ro��E�0�#na4f���j)���	zU����^=ԟ]��@�dl*c����!�L�h�N��x�|��^c������d;�@b9��z��wͯ/��UeV���Q\(�S'�����D'nĠ���+D�e:�{���Gcڍ�Ϊ����T��	y��/q������HT�����B�J ;x�����zD"�*��	n��:oI��T�Ȫ�9����Ǥ�
Ef�'���K˓T�64�����[H�b9��Zا�su�^*��^����T�w}@��.�F�Yh��횰�A��4��:�)?��e����.ɔ�c�~*Ʌ����3�	�ʨ����d=#��G^T
�m�!T�}�kYe�w9�i|x�1K��
�BDhcD*g=P������Lȃ*�[���k��y1һ�������ה�;rv�p�-Ȉ�n�r����/`{���@�#Ĭ�S��3r�	�K[�B�	�n�@�ӱ@qv����{�<0oOe6���z6��F�x`҉� ;#�'�����j�a�ILa���~X9�_/���KA��1����}ܿ�g�q���=!�	�O�2:�e��������6��g�r���:�q�ެ~1"�<�'s�O�o���^%��)��g�=�3괷<�xC�����P3�h�r���2��������ZCU�{5��?N�P�yj�F��w K��9��E=�0�H>��7�q�{m0|��y�㴅I�`螱���4��\~~}�?�a��C�#G��{�ԧ����q��wn8w(�uC.�%FU���*�����ר�T��R���=F�'PM]��ɭ9�	ɴ2����a�"�_������ˣ�~6��W8\�,'�\4�k}�9�7c
5$t���4���S�Z#ز���<0ڌvl'>>�r^�y���{�����n3��M3�$�S��,���or����	 ��Ω�b��Q��5ҧ�;#���u�WY�s���$�_����a�׼ڿ�N����>�"��?�j�c��=������V�$'g:;ҁ��F�n��h�_\��o='������&�[���ˀ�[��a����������c$�����t��2�Lw���g���=G���
�l����+wA��jd��I̹47���r�py��!�*�>�5.#�Lӂ1ї��Y6̾�V<���^I4��-�]�9m֊���[#��c���ҭ�z���r�jn/����*�aI9�ׯ.X���q:�=�-0f��f{��c*�a�Bk����p�R�@�1�`|��~hQ�-���cA�
|����P���G����<�ozYI���o�H�Y��X�	:(�J%���U�Pj(���AV`��u<�~I��z�U�q��[ϒ�m0;7�[�y�)����l�^{��"B7����U�H�+���-k�y����!q���F���2�݀Nd���Ef���_>.XkD1��;G���[��S�x2�G�
�b�v@8!���%���iR+��Sc�3/�l�o�@��_�-�&)��s+����Ŋ+HV�挭��s^f��9И�_�|������е�.�0w\�D���6a7t�|������!�>�0?�8�. �k��םg=�!���h�a\ӷ}�y��M�(6z���>�\"`�m��K�r�%�$_-�T����3��;A ������Y:d��3��	;'nt�4�S�Џ�x%�L��$�]pD����+*p�+�s����%�rp৲�u�7�W ���\�=}pk1'��kq�G�pd����<?���tʁ߀�\S$'6(�����<���f�<��̽�܎zQi�<:<g���59ÕA�l�_�j��S']éarWu��C� �G컑֚
��Ko��^-�:�w��A�׺�^!�c>�;�6r+0�1�ɠ��4NM�5W������|(��Z��n!a�B�>i����[-�_w���G���C�BAB�:��L����EX�n��?�F����-�;��L�W����?��H����8)9�P�{��-�������S�f��{E#?(��w>��0l}�l�^��h�)�?c瓷�O��^���Ɲ�����N���2
k�$�mI;�%��tw=��Hi� #�n��Ŷ��ۮ�jM1�ы�5mT���/�12 ~>��H~b��� � s�UȡMڥ��3-�'�D���V/�g�^p7��l
�!�A�ੱ�!��5�ﱮq�1���b����J�TH�p�
H��)�,y3] ;q/��S���������D��r��碛%��m i-f�7��uzq�%�������/�R�7,KJ%ӯ2����O(��n� 9�W�GE�E���.�$��}��+�.�|_�a��%myct�Vߤu���/h�B^�gNt��,*hw�\[���0�5��i�+��J�R�����ı'7c� ]��ܤ�a��ʬzU�w|�~,VY� r�ڻTd$M��fq�кC%��!�Z�D��n�xs���G���/����-��m
{�V�d��r!l�=�5�
v�P��ۈ�C�X���� ��v ?�m��ߗ���Lţv�O�ޖ�R�(�J6!ڼ{!7��DPXI�ݶ'&V�������vS��1��R����Q���� �3�k��:{_UF̢!ʙ��'�=[�A�� %+6w{��������%���s��	g��f
v�e�y�Z΅���0�&������7y`[�Ӫ�9E��|WU�݁+g���>vM'�� ��jߝ�!��rR3�#)��g���~����5W9yB�d�sBnz���J!��n�5���=�w�YĊ�����ga���o!�vrk;E�:ʵ�p�����T����$���'���	�$����� �M�Q��s�i����h����*�(㻜��~���;�b�c��N���oUzє�6+�C���7��;�dؤ�-vm�SDc�C9�m�yME�4�)=���Ţԥ�r������BC�@l��V�m�Ꮿ���5O�q�ָ׬)z9�jl~�0~O�܎n�ą�m����	��B2\k����G���c8���H�^*EgU >mSIȍ�ܒ
�F��JrfF�aL��ˡ_�7�H��A7���� b�^�"�G��_�k秓@q�VBA�~L�&������o�'9���\$}\,h�)�&u�s���={� <{�Tbޣ�}�wg׍�m��2�D(��a����Ύ��g��5_3�Wo�Ж�o�X��W	��پ�	�l����}8!@	�D�!���ܡF����
���^KԼ��I r�a�_�+�9y���U#����(�V����ힳ�<����Tq�=�/�a,i�4��'YS$�I_�K�-H�nk=�մ�����Kd"���A�I�]�I#�x\p4�arG�Y�BH���(�*�K�����a)���`����kJV����Q?P��I��w�����>�:��\��1c���.L9D�˞�5`�E��|�Z ̈��V|
�*,�bQ{�^�1�X���pC�^SR�P�?C�KH�9t��E�O�Gw7�7��7�e�/�W��X�S�T;ƹcZ�9���ힿ�f��4nQ�G�m���Z�����;�l6�w�w�Hovr4�7s�k�Ie�X0	��+�)���n�^?h<w�w���"��k�-��V��᫁�>�U���/yJt�Tf']Q�K�����J�z��KL;�ab�E�Ii��$�k�a���[���G�ۓ2��A�B��h+��pmX���:�>�4,4X�OW]�|�'�A��Yx�w%./sZ>�O���瘿����Ob8�1�I�Ք���a6�bk��m�G��Ao�� �bnY������h�� ������ 9��Q�,�xq�h�z�y����Z'�]�.Rb�",t�6h~~�!�ʓ�W`"I;5���>%u���������hz!�x�,N�6H�8���7Z�^6���ib�Lx���/k-=H	A� n��upLo�)��|�K��j�����Y�`(x�$���2oELj��=��ܳ��c���΄2�.��-��k�
-*}j�L ��Ni�
�^`��ƣ�&w+Am�x�MI�}U.p��%�Z,�6<fJ*���uz��v�B�*�xL�.D�4��`s���S2c�z�m/�h�Imܳ���-���7"Ǡ�U�p���&,9��u;8!q��~���A��r,]C<ih_ ����Ն���D�7�FJ�=}���&ؑA��/�\`�[+�uS�^�2��J��s�e��$��UL��΂������`��
4��:�'�?�?ҝmQC>9��Z���ܻ���`�q���ה|�vQ�2��8o����D�r�����,�?5C<�ڔ��A>r���D�`��b��nc��b��]}��*<U��V���Qф���q���O^^���7�����*�7�|�«�o�&Z���,�r?zϻ�S��Ɩ��ѓI���|����"������XM������l/H׋2V,޿�p����	���{#�<�87�b�4S�N/z�|�F7�f�:����PQ=S�YK8 L���ݎ�2[走�ʍ%Tz5j�Mw�u����!U��_5$N��n�G��qB1� >G�B��Ԝ�	���B�n��/ʉ�U�/Oqv$\�:���^��i�'�4�S~��5ǰ�Oi`5��0	�k���v'����Z��d��ξ��-���Q�1���y�Q��+�������0L%�)T�:���J*%�~`�f��k���F�2������,��#�b���S%�`�+ ��_�b��@�)��P4r�[8j{}����48���!��s�m���}�nMbU���}�cN�F�+����Y�tv�O���2���V��_�U����lx���l����g� Oɐ1��,�&HH���_{�\7�?�5c�����'�i��	�Z9�ߵ[���ج�
����ZdD��q�ީ�ܧG���/�Z5�#T��ObTz�Z���8�%�f8v�����b���ZQn�{��&�����섪��Qt*?<Ҫ��J-eQzn4���Cc��V�1�{7i|�h������%Y��/���\S�v 	�]�6�ħ�*`Ư+��1ڬV�xp�M���=vr�e$��?��ht�ty�_�ۙi�"�E�-p!Hq��y�!���9��s#~��苢�G���\;�0gR�~�f�Z`�AZ�$=�����&ܘ����fp�ޜ��Z��g$���7+��J�)��~M���}��q
|%�Y+�N�/�9��a�������N�M�:��z8�Ⱥ���"h�#�� ��%0jR���e��  fq��\�����#;)n����J��������1�2p����O��f.�����>��v�+BY��y���	���zvMc'��as��UA�v��+r-�)]��ӌ<��vt͍��/�U�������n�"���x�(��\�$W�@�pa��B u��U�w���m�ݹ�YQ��ez_%j�/���v�Z����::�.6h��O��V�P���	�*3��;�@�n�7���q���u6�]nI ���l"���@�ɳ��)�
�0�%ޮu+dFiP�l��n!�@֜3/�>����0�����E���JF�A@�����?�˙���*��dc�E��<"��@�!)K�ӧ�h�;�xח5�ۈ[����|��R�'���|T#�`��`��(x�eK�� �1���_JˣIANE�w� ��(hHr���E�ک��?K��$�F��
99�Ϙ��$�P�jx�x���*Q�6S3�,~Nj�e��{�P'[S����3���M�����Yg��W�(V�|�{"U�JV� 
�P4���(BY��Cu8P����r�+�*�'�-Cu$��L��\��:�V���޽�M�_lM�jʗ�zXe:Ch�eѐ�5���\	���/���%�/�msX��m�c�����ј��da��b�6\2X�`�X�i<H���nUի9����1X���W`$n��%A#�APIa�>x��@<3K<2��M��\����W�r1潀<�3��+6"��wj/���������f�SG$��}��A�%�J�
�u���`�	[=U�s
��A;G�|�wz&G�������@g��X��enBw�E��Οj|�^E�|��YۨV��/{��W�,��]f5�ڔ�Tp;�c�h3��3�g�U�v�Hd�Ț�%�����d�k�zF��r�z6V��81w/���sV�-�{Q)��nТC�5������ă�9˩!�MRU�y
{q��U�������#]̑���s�S���x|s�Ƽ����]���8o��-�핳Z�{r��N����QA<�D�8��|���o��D�.���CF%��|�ŖæD�t򔸄24��"<�Ld��Ѩ���v��Z��GT������Ц�逩!��� B����o�۶����+����-Z���L���&Ô�����F�m7x,F���&�OS���˨��v����\y2Rt���_ϳ�h,r�P��x88����À'p��;�=Ǖ���d�s��˲�j�;Kj`�Ǎ8~���}8w�$7�Ыâ{�̓Y�-u�BP��:�=f PZ`�f�$�J!Z5���YXS���W��2��B�����O����$��&?�Ht;�*�x�2�M�����%�
��"�Vׁ@T߭06IKV �d�7}�6D������2ٴ��5��Su$�1��e�A33���t+��u����#U@b���R9���~�贁Λ*���n���RW�3+T`f������+����b]�'�jp�G��BP�%薆]T:���"��U]!ˏѹ6ʃO�TKB�Ƣ�D�#�60�z
����rz��!b�ר}��,\��G�i-��+Ģ��D���=
BM�jr����LZ�$�����&�P����0�'�jdrԁ\ױ]���"��P_q޵�2�������C|E*��2����n,������ߢGaNț~Q���;�zH�z��A؋l�'ސ���PKv` %�-8���5��D�#��b*�&����C����ˇY2�y#�pA|��I��1�F��;���O�b���;D�htؕ�����=Hy��N*G$w���v�zg�; P+���j{	dK
�k�/��.R��
�"k 	��@X�ۋQ3�KPG5�:D���� y�"�O��W�4g]j�ނ��vt�&�>6	����Ы���$���##R$� Se�J$Y�e�f�����wX��G?�V��H�z`u]�,|O'w���B�]	�d'L���|�Q��LN� v����Zq��֏���I�
��0-`��:��m<��%8N��	�#�Kh�DS�E��U�|%?1�ϋ���!b7 �Ugƛ�u4�h�xzB��'`'�<�\�����x��nx]FhIT��d'ј��o���,0ήE fx��Z;m�:�P3�=��G���P ��������[M�<�Ĕu����ZrId'k��F!Tre]��j��|��5���9�=I�N̫�^g�v�D��zv
&_�I
K����^�r�!�ÿOkt�I�K��T�Қ�r���}Q�` �/��I�8z�2��.h�˱�i�ٲQ�e�n��2��	W�Ō���`�n�~�o/Ӣ �D�t�e���Yx`�@[�zB�e�̯�uMo��7�%6�͟�2�02O�78mu�Ls�:Y1�h�A����fr�Q�d:���yt��x���>}t"6��ՏD��ǒ�KΨF������`�.��Ѯ�4�@��	��XӰ��:�c����m2���Z��euN�ܣ�i ^{����7kq{���C	0=f�]�c�|2�dWiB�E��c�bK����AEy�
6�L�@�����ll)S��
ɲ633y��6�NG�W�9<�	5�>���'�[����`~J#nþu�Mpb���助4�������{�<D�[��������Nŭ�p�=Ƀ�r�߳��-�5��:QZ��I�e�`!�y�+�eھ��/�T�4��kR�I��\�Lz_֩�����qG���4�B9���z	�ꍃ�tq�T\�|�<�6��m��~IcL����밨v��Xz�b�ݿ}�T�w��X��`!º.�w��{��Uu.I��Q�����1�s�^���_хT|�Ʋ���j7-#�����z}o�հe
�.j���J�T��O�jB�R8]��[�	������>Yc/r�{�&�
�k��>�ۥz�@R�b�Y���-Ec���6�6�^���mH�0H৆�ؽ�u��k�j�G�?���a�lOP���!�i��ZgW�^�*p!�T,�"(˯nx��9k*��V�;���+���N��3��xD�"��ŕZ�1�ք��v8z*��CG�#sy� ��+�f�Y'�m�9i5�њ��o������Y��D
UNH�Q�,���sR.���W�H��p����T��t���R8�}k��Z#Ǣ�1�/)���f�^4�I�E��>Lo��f�٧������b���g��K�����.�]s��AL��q�FS
:�W�4��ixh9K#����$�V�~� �L�v�������yo�~YBkӈVM�>�m��=.h�v�N�t��ֲ�&գ=�[��u�U��1
�)Po;����4�!�����s̲�2<�v}��/�XU3���l��Ǭ��тx�_��A}��5��8ུJn�޿�A��  ����cGag�p��f�%y]�O��ݴ� �4���.8����dW�r�4���g�H�S4�9��x{'k���Ʃ����3��l�N�ҷ�
�"a�B�e��U/XD�|p0�l�o�>��'ڗ(��%�shPj�sSe�8���Q�i��g��+�k@o��y�M�c5�vۈ���x�)c���IJ�ĸT�H�?�K�
��B�jC��>�?�����
�؂�B�+I
���C����vdW��	L&�˟��^i���L����ir���_�Qv�I_�	C��p0�]Lh��i�������X:2O��3f��ٻ8�!Xqr)H�UO�ű��FPU�+�6�����0'l�v��E�y���d� z�A$%�xK��=l��Mq�CQ"���i`ü*zk
�x�k�YG`'YG�}1*��U���"6����[D������RZ��#x��|׺�`
�xD�-.c2�س�CXÞ�pI���O�B�`|�Ĭ �HZ�D���uScyy�m�xF[q���Ah���W�+�AYe��M�Ac�i�&s�b݂^Y�6;�}�:Y-D�`w^��m��^Z%�󌗲�/R�,t��@^z�J<�k4�X�T_9�$X��o��V���a�4���ȍ��|o��"ok�{t~����P�lX=����bE�7Ձ����H���W��w��ѡ��7������;t��u�n={l�2��v
�j�:��v�,Z�}H��3���I}3��\��H���
�ö����~�!M,Bʔ�x���J�^�W}�<�z�.�h���m�M���i�kXYS���`o%�#՝��kv�\��Ku�TpG�1�/���{ST�5����F��,��~ղ bѴI�9�e,����{�&G���&��J��5�!9E��W���6:t �hT4M����C�`����yT�����RuרH�J˶��J`%�8�RR�j|���J�����7�tB�L����NSS��%���qqT�[{����A �D���Һ#j�Ǵq���#rhEn��=w���H��0�'䶿$}/�fT�Ɨ���o"$���ٚ��lŤJ�
�����ܯftFнٵ�s/v��1��}R�+��[��)2EqN0�e�ۛHv=��w����Ϛ�.�U0�@*-���ġZ��Ȩ�u��,ҽ!�0eg(_}��ۏ�3�m�y�v�}�XS/���%.��_≙H����9�v6� �t4ʿ���R��Npr~�y�l����'��ƬR�?\}]������k꒎�aц�����Eb��6& 1+&�~+��@�1S�<B�+��Of�oO�~BR�f�)(����[��3�����L�R4�5 �(�e��[!<Td�3���)�s�E,5�E�tY���^�X5=��K��fU$��n���,��5 ��M��v�r��w*��䰟BJ��K}7B�Fǲ�s�G���_��X�1*�ٛ���&��GR��A�I���I����9�{�'1�sZ�KOn���rѢ�pK��(F��^�\�(<\���T��j�J��䘑XŰ����TF�4��j<�zA��o8�|>���u(~w���u/T���h�v\,��ֻ�w�s���`�C��lcKԧ3'����\)���&ŝ�f�ƥ��Y��*����):���]t�rÉOڡ�Y<>�)t_H��˿������H�|!O1�C��x��s���M�G�Ҏ@q8�p�?I����7�ic��E Pu�%LJ̡�W;��qF|1������s�VnP�$��6�&!���v�dg�̑4|����N�mu�*Q�q��qK.8+�ȴE�S��2�q
|O�ӏ���P��]p_�g�@�e��E1��,�c�u�U�9=3��b�S��@����0܀�_ܭ�> 	;wl��t����"���AM��u��e��,D�$�De]��%�馼d��p�NS|H9F=�%α?;<��`��u��I1�����W��rw�'��'�� ��mZL$��F�f��[���!u5�fԽ���`5�ƌ\�a�-���z^!��@�G��В^�a���|,���OĬ��,z�C��ק@6'�����r�C7s�n*���wy+]�E��RV�`���E�.t(��>���rɽ��lp\zȫ�<������;��1��K�rP�b� �[��Ș.d �z,���\2�g��9��}�k�M�$)���D|���0����5G�.���!)�juӡ�c�Pu������K
F���XJ�Qx,4p4;� B�D�ܮ&uk�D>��][����h�R����<B31��n��MJ�4���`�V��������4z*��:�'R���r��ߡY�:���Q���6<FF�"XjN���LZ5�в@�����^��k�ί4���4��ݸ�u�+4l�k/���W�1HMȎ��|_�f
 nR5V=`����AA&�v��aJ.r`�Y�Y��Q�X���>��/�9��Q��j�\�Jߞ#����Z�'8�q�k��Q�,�
;� 7V"�"1@_O%�S���x��00���Nˆ�QQ��-x�i�AO�J���]���ث3�#�Hc�X��"�G0ґO����Y���PG��J�H��^�g�7&V"e��J;'Z�ֱCd-�R�X�\���8��b3�@���덆����!��-4��������S�f��l�3�L\301��U�����H2DO�}���W��It��/k-_�Np�k�n��G7��Vn��<��q���)/zQڑva(������iE|�i����v+�j��6��E��P�^[�����M3V1\����L/��G~���7�Qa��A�Ghtnqo)d[4Y�Ob���d���Pb�NN�~��P�0��	�ULt�ϩ�wA,����T�7������>���y��%��r�,��o\�?߾�UK\^_+��k�[� �j��s[���� ���ӭ4?�@�q����G��)4�½��?7�DL;�6�:��_�H[�9���vcx��k5a���oHjJ�YM�nfZvL��Ο�DX� �� j���jpIL�x�R��2�K��f =����2c���������5#=~/?��v<�hTKz\�\v2O��a�(�5Jw>�jW����h��x\R�-*A?"�r��| �41�^��_�uYHϙw�PJ�כ���\;���jQi5?�
���ZRc1����oz���6��iG����N;����k�8��^�I��?�/�GVm�|�-���� ��85�P��3g�6
6a��p��*+x���%Cb��*����9�I7���`���'#呧>����*'��f��A�~��q�f읤W:�ǢXVR �һ~gC�k�̟�r8���t�xW�e�
sb�����+vj[Ұ��Vv�>��_��eݩ!ݸ�
fK�{�w���	�ɚ5UX�����VZV�!E|�#�f��.�<����IEi�D��0��*��%��nRQMP<�Te�L�@����)9�ԙo䎯$햰l.��Pu���+�h�}�՘3��p&��N�����Lpr������F��G��Z����	��on�2���6��G0Gl�E���^�J���.c^٬�}�~ã�V�ԾxZ�f�dA�x����ml��<M%or�ps�������ok��s�.t�P����o��rrO�,ԇ�w�����Q���v�f
��F�\��M��(�t������J;H���X�+R���I��=<��Nib��[E�5�j���� �t��Bo�X�(�b���O=��7|4,_PV;���P�̾���E}B�rc���kwGE䐉g�O��d��u#���I����'WQ�:�4҃x&�r{�op��0�2�}p��1��3�q-�4[V�k�@��;G�5��WG( -�9Fk��
���6&�����d�xfzSz%"�1|v��TQ�N�U�l�"����^*���2��FQ���|���E�0�����K<�eb��<������#���.��Q5=�$�	�B�^�d��Jٴ98!g?�힠�u��_���9�G1Ǡ�+! ��p����to[^'֖^�԰�W�++}jE�����*���&j6�V�/�ƃ��k!"̕4*o��v r��T��\}�ߗ�Z����_��FikJ��^򱗓C�l��d������@�BY�?	��8�"*�=��g��?�����p��L��'-�l����;jHS����Y��׭�f���a��{��z�GjIGB����Jb���Bx�
��c�~*o�����/�S��Da�D?�~w�C�V�IG�c��6�T.Bʃ�z،��ً�Аn
Rf!bT�V�WV�%�i�H����>��_�"n�B��:u�k1n�������1�D��QbV���W����E�C��-����{/��r�vF ���O�CtM�=[k!�	�7�*Vi�>�h������?������A����u��hЈ�}-w8�!�f�� ���a���x����4�e<?:{��o�s��1&�e ���b����I�o�X����{yx��s��)�¦���6]O�K"G?�ӆ��%���n�7o�iѹms�Zo]&q1�s}��i)�݅4[���e}Ѯ��7A&ErCd�ԃ����D�
���HV>`q+���$��	G"ȒLY3�^� +V���xIyW�93
��ZVg��S������g�ZG�:���L�ݟ���1�p^��=O�П.�?'�c	�Hc��A����G좷�LADRHAL�T�O�f��¶+Z�M�̚8J_*Sh/���d��_��R�cبm؉~�;�[AR�C$A�ټ�ys�+��PU��ߒ���1��<r���?���&�j:H~��"�U�ۑa�Bݭh��\������NT��y��gՉ���0d����n�[v��󸆐�"�6������P߻�\}�6�_c���S� f_�R�tD{�@�e���Q�J�Yjl�e��Es��a��5���a�m�Bg���z?'���H`�����w�]�f���J�+�p1gp%(��#_��&�N-jI�R.q��ھ��[d��� L���$G�����$�ђ\�rw|/hYC�:�(�W����v�<�{(�S�\s��N41Ѷ�行��gI�*��o�`���"y��e�?g
��(UX��Pr��GK�8G?ݜ]���7z酭+yOJ�l�ތ����i=I�3lw&;�� ��Gm^fF�� *ω��W?����Wn09��,��
���\1{�}�מ�lI�&�����mU�|�ں˼?�p���vx�lKWk��*9�fn�����5c̚�&�)�H5��~��Ҿ�M
�(�ݫ�1k���v��0~� ��YƔkVTұ�5��!B1���g�Wf�X�_�J�]��
�tD���H�#m�%wi���iK;�юhEʦ���$���aO9� �֞�i	ܐe9mDy��]�������,���c��A���x�,����N}��~LM�т�N��
�rww`���U�b�kz�s���Li�߮���o�%O�6{*�s��2 �.\�=�C��em���	�ӀClo���շ	�I�^�]^.��ϝhs��L��� .a�G��&�אx��h�b�����wI�57�FO��ޢF��P�)�(�?[o�P���/�߰j�Y�,��o�s�1>�st�CI'OO����n�MQ���(�$��V��ςX��X��]�OfJ����>�Xib��J��f�*\�v��Mʻ�o�|�9�`��U70���y}"��>L�@�X\q���W�_�	-�!�TБ�ŲA]��Vi�����[K,�:6��Lf�j�L���x��NY��bU-��1<c����&�]���qȕ��V�zP�j�L���0UT�y�	�ؾ�Dɦ��W��Ղ(��2eV��SK�E����V�8����0HKo�����v�R"xX����H��=i��5rý�c�%�>jPEH�s��p�a��R;��G�9^���iË!��G��
GJ�7�E����,����ۡ��K7y����5�"L����,J�}P%��W�ֺ�\����c_�r<��!��GbH��mɬ�I	\N ��P���FQ �r>]�yX�<{��Q��9���#��v�V~m�)���|ǻ��p��̀�1��i�l�����3�����Y���WT�Sl�|@$9��	l#�g����O��,�t1'�I�p<`���띤 ���<@'Sj͕̊څ�)/xn3�Z�%�O;�,���&��Q�>���8�s�xg?\uA�6l��h��h�ס~D7�p3n~%]Nd`�[�i�^~(D�*n=	�e?���!R5!��[�ܟ� ���+�E!sm�7r
f�K#
�=�m\��i��Z��������L�U��P読�D�9U�!�PFm��#���&)7 ��Ci��.����,pSD،~�=ߥ�JZ�ш�e�l��5�N���2�<O4M��7�a�ϋa�ݰy[��]�E~k�C��E��a4N��>H�Q�4�iULeYQD�?YHɬ#�y=l�C���p�I� zV�6�_r���.⪚7���Q���N�b�t�ȝ�F*ɖ��s��̝�����^��G2C��9�U��8�pݒ�����7k��E\��ن�i4c
rLe��_@Tg`)\�_}{.d���o�w�� ߱P
!\�d?����]�:���y2���4j�Q�x�:�$�E��Y���\�"����II	X�Ae5Z��i�J �ٷ��;�Ҩ�ꉖm��]$J
O#M�f*h5W��?��>���H=���X�%�Y�h�ʹ�0��/Ш�2\�J~M������5��N�鸛��e�.��1�Q�֭���k��/��+�S8iՆ���#�N�&��� xhq
xLЉ�O܆��b��!L~���p茗�<9�S)J�vJu@n�V��K0L@�ǜ���E;��:{:		G[^ē��%ǿj�\�W�9���:�c9T��U�2�٬|�(hlTj�������P�� ֣�y�c��q���1*��s��a���k94��Ovb��_��.>�����F& *�j�����𠁴��=I�C����RO0�"�V[ ����cPYm�C������W�8 v���h��4�&�Iw�5�t]���4
����k&�<��p��% [Q ��ƒ3D-���0o�t<���I��v�t�O;M�8������֙i�T���e���ODB��z"����t�
�ӽ��$(�k�'CsF���I?��W��cq!m-z�_ʗqw�c���t*���c�wr73��W�	x^]͙�嶠wW�7N0"~,���aC:?�e�����2��E�:������&Ii�E��@y�H5��7<�!o8�����.����{�\=�i��B��v���r���x40nY�?r�bۧ�-�dj���h���_���g��wq�Z$���?4��x�r	�Uv��λ��������ncYZ��fYv�����������.�>v�I���V�o8j3�m7&� �L-��X��<RRB�����K�¼���B�Z�����Mo�O������S�,6����z.��)d���F����&��$����^�g?��JD10<����� �C�gP-!ęBoX����b�<�	�VR,�1���2��P���~���F�M���P��	�y����yQ�<�vb5�����x�$���V�3�o*}y����^�����t0P��?Z��.d��oL��0�Ґh��l:���	�������Zz��SIXP��rL^+��Bt�A�+5��Њe+�f��m�ӄBL�M���z����0B�)p�K��#��vV�n*�4����ؙ$.iH�'m?y�z�����Wi��aX�ݻ��Oso�"ɕ�? ��2�-�7�c��r?��8�9�v��,E,��M��������ɌL�6b�v�_��o:�ӕ�ފeBe��0Lj����.`���#��;��X9����B6Ʈd�̥�T��F�:vֿ��md��Ĵ�"�����t!�~���18W�(��JI���v�7X�W�`�3L�g�`>���$�1�֜WF�gL�@�������D��Y�	�����?ި�,TuJ�n��_'�@�G؝��,e�a�4�h���$+�?t�Y<Sϟ����6���eR`�H�k���z���D�.�uy����D����!�H�8T_�S����*���Z%A�/�!R9�9���]4>d��E�U?cO}�*����e�	���)S��/B��nj�hg���D㱹��!��H'��e�ER�-���U�(|N
�[q��f^|��J�$��U	�;N$�L�a� H��Sސ� E�ٗ+�	5����9��n|��^� �7 �O	���u�ֱ��m�l^5��0��P��2���ۥ����ţr`��t����}R� ��;��^��!��Ay�}RV�h��L��\�����^?h���$�����Q�d 9���ʴ2b,�A��l��6]�"r^c�D`:dF�U���	�����>��X�Щ�o�/��<e����xx��RfI�(�)�'ո�ŏ5A#k7r9^'�&�<R*{������v(>7�џ\�m�o|)�-�����V�|�Љ� ؛�֛�Z�/�5��.�O��@u�z=������6�vP��j��K���8b:��
S���Z���(��azs�3�1��"���C/��c�η���T�u3W_�V�=
�Lx���v�$U�V�x��qw_�$�F8�K�;�mh�p���J3�R�=�y3���f�ߩ�E����>�S
	no��#�B;s����ūE۩YC�u	v�Y0>��Sn`Ps�pN˷��#z�Ak���Ñ�E�����D
h+�]$H8�㑋�ql���z�>��v��~Ú��d�<|+p�Ǎ~�M�5�)6��'��Q&�d�mz5��Ƭ�#A)�Lf�ƁE;`�i�3t(c�1��gw�c���N�Y���+����{��Xxl��t���yO�2뿨� 
�-]��)�5/͘>��∺�;5�b�m �w�G�)��/(���MI[�F9����R����=�2� O��%�E'Ze[��-�p�w��q�n��]#�B�tR��1���,L^���%���$F��;�&���ݣc�jUS$�ql�3�C܍���9?A�z�~d��qkiJ��4t�Z�
R0����W�t�sD_�v����Akه�:�/���������������g�{r��MIC��J�͝/��vI���-	^���iP�m��@o}�L��+�	-.��ᡜ��l�v���Y�H��3N�
�(F*�{�Y�7S��|y�z�{��������s4��'u��n�n������,4,�=�˺ݗa�;�-�m���Yy�;ủP0rB�� *�����4����l	��6��o��u�Rt��p5�����npP+��3�'w���
��#�Q���� zPJ��~�aF|b��27>��O�wҹ�8�V?:1��hs'[�}���EDv������������`+Q�n���Zn`v,�T�ϝ�L����l��Z���6er�b����e<*�� ��n�����ə"��9Q�R8hkܞOE�-07�us���ӯBw�Ή����2 tz>������m-6+F�5c�F�k���j��(�9�S�򚤜Q��*^i�Y)�}�3!��k{�a�N�e�c���]֔�I�GBUc}
`��s=T35��&�ֆheo��*pU嗏�S0�l����9��q��]�n�5����1T��"��x͋�BG8`�W��z��M�-$��P�K�:Ұov%۴���$4`�����s�!��D�W��w6�7�nL���Vs�&��[W H��r{��S�ܜ��w���G�m��/B,�5���x�+J:1w[!+�HD�E�f� �w��6x�0��g./o�̅qaFK�ֵs�8ϓ)�8_z$���5�3喊��ʢ�/�!J͈��+��)���O�Bʇ�-oN�A �*��gH$-�bKw1}4������ܾ�P�y�DѧE��@~� Z��:�~gBG,�y}��L�c �'�1�-�z��"\�ZOxCa�Q= ��*���g����p�#�٘���'���9�qi�A��(^��b�L�f0n�ö���h�ڕƩ�s|f|3%F�zK^��OY[)r9'�T)����V�xv�0��ܒቿ{@���s�">y5'J
8����?Y�!�%}ș�μ7",E�?��R��j�U�h��H��G��ZppX�<�9F�UT^x��:�RPh�2�AW��;?~��*+�B�E��x���oD5���F	��
SE:w���`N0��G%�N7!�6nr�_D\վO֬Ձ�l��8�U.��J6}���A�~eϪja��\t����JQ���	��ɷ�(��⚣���ù��w�|rӪc6)O�(�e��;�p�Y6'C1%s��M�v)�I�Tpz��].i��Z��
��-^7r�^UT���q�:���+-.�e�q?�++R)g����u $o龅�+ћ�Y�_���NN�������机�G9>������C(o�ԑ@�t�b��	����6?v/" &�(�&�phF����������������a���/hIc�sK�a�,�ʪ�|5�gXa��(����EW����y��K����\k����S�߁����3��Npwk�RI��S	�*�/�dD�@�X��L��$�'|�����ã}��\���T�Pb*4�W��i�ڹ9a1t>=�\�%{V��}�0�� e�t_�V�jN���歴��i�<+����7:�Q���J���uf9� �1��A��:cO��-�b��?PY.%�������I0���Skx#��(��x��ڦj{� E���r/�h�cȖ��"Lco�Y�A?^�3�ł����iڂ8�>)I�^���O� �W}GZ����
:0 �]4���͐�a�s�v��_^��k��ㆂ�Y��%�s��>�@��fx����(v��I��A��F�hF�~b�d3y����5�۫D��A���o�Jl]�u{���.���h ]�N��z���2�s���D�}u9ڈ�_�H�I���'�����m<.��g1Mf9���(p!���&���Nk4�~�ղC��BM���xt�ntIE�g'��y�J�5f�a���3ݺLtط�_���5�&�G���a�����Y�����>�+$S�9`D���`�pߝe�F���S�:%/�`�G�Ђ���VR%���i���8����`��F���������G�R?���م���	`�2�0��R0�����z7��b�5	r�Z����1:�iİ�|�>�~<�æ^]���QNv[�M7�K���4 ���4q\������uq�ʫs�npF`� JJ�5���;��6[�ݙ�uAq:u��JDmmȦ����2���畄�(���H?G�ϛ�����2Ajɡ\��Q��Ou �n�)$�ˍA������W�����Q�e&�_2D-n��aK]	"�E�y}s5E .Ĳ�U��aP�\�{�D*:,]���8��y�����|4�,�*5~GW����1���7%/�F�
��%k��Z	p�10K	�6�.È/���H�Fe&�=�����2��|/�EA�;�����������L���aƢPz����E�@QrN���%���*S��z������+>,�]HNX�����jb݁��Ih5Bpz��B�K��0K��J���/�F�H.�_=�с���`���s��XY[�M�Ǝ����c����D
×����@��Z�Υ��$����ӔP�)�uu�S��/��X?���Rߏ;����xp������6������-�d�M��j{N��Ss�ݎ���s<o�5j���n��_�b��6�A�X�G�+�����9�#�6�+
�p<�^��D�Z&�.��*W�mV���b���/�Ļ�6�JB��/�	�dɀ�a�q������E�Ug`̡b�N� �;׶- ��sc@k����V��V1J(�2nt1�0�ODʺ��7o
�I���������c�"��*e�};��>�	v�=]��{t��e��VxS�=y��$�r��9������Y�����4�|w�[u���]q��Π��D"���q�>`ɛ�P>�^]ה�!Wj+�q)[�t�z�7��-�}�/�Ť���t<�g�%���Jʡg�i���?�߮�U~c�`�@��:�ě�d�ۊC{��u"���/5�T޽����8_��+jR���`���"�@w<m M^=?�S���l\�x�ϴ��y띋��R|�у�����m��݊h���\�c�M���6�Kux�	�5$s5�C���6���B$�ɑE(d�.�^F��� ���
�/]-]��پ!ʘ.Ukx*�	���Y���U��y]�dK_�+���GQ��#���1��?����.����<ajqc���୊����4XT�ͱh��ix�OB������>�T�!��֬����/G+!+�\F�HO�:})����.�)-a�,���]H)�|�s�����m�_��F
ڐ�����CpPhE�?�SB�ėG�>������|�YQ�8��u.d��6<��\�^�)��/c��_?����g���
Z��*����F��ʌ�s��'
�A� _ ��%�*�
�e��k���8�/���ߏ�N�`�9�EU�� R"FZ:��m-.���7t,�a�Z�Ym�+Ǝ�'���{*Q`Y韵�U8�@(Lf��UK/*�x\q�p�d��_;<.�s�ݭ��.A}f�?��K��l����3���%�w�*��jy���J��IR@��Jg��fw���"4�+|h;�TR٢��D2�ћ���M�3���tr>�0��F�硇���A	a(�/���D��?��mRP|.C,��[�t$��Q�j�F�E
�z������sb�O%��U�y+���I�U�Y��A�%]e�`U����-�(jX/0	���o+M�+� �m�땩�6���k��[K��:!������h^�}������Qh�����ׇ���,~��'� ��M%�`��p��9�O�L��0��	3��o~E�_�`c}Y�8��B*S{�\����[/� 1K�3�(��$d����~pSA���������N���fˑ�?ܞϟ���l��;�/M7kh�:�����x�DM�)�3-���� #��J�1R\/�.O���~�������B|G��z�/iЎ]�({�ƛ�D�שz�X?�Gfr��S�K?���fx�(���S��z�d?�{rI<����HK���5z��$���Z�>�.+~>�#�}���A�m6be��L֊��������:�?p����X.k����(9�F�W+D�u��i,��`7g/�nE�[�2��R$�.�C='L��rL��q���g*��:�����@�����>'�Ď�����)��b���!��)e�X��1���ɲ��WQ���\�hBm��8o�Mi"Յ�����KU�]6����US� Ųz`��@[puuȥ*��>]�V U�_��G�u�J�>���%K�~��M�%wA�z���s9k���b�Zt�v�?p��dpM�7HHpmb�� �.ޱ�� � ��N��>7OJ�����.�~� ��֠�HX�GS�'���r~$�0���(�ъ~�[�)�ͫI
����9V�:�C���WJ��Bu�X+����$�[~N2>g�\v�h�D�V�i3�e��޻���3�Fܸ���U*�p{Υ��.-������L����Ie{��*��*?)K�+�>�X��Q��`Z������������3q�*>�����
�Z��o!���E�%�
YX�CNHc�6?�%L�z'�=T��^U;�V-�r\L({��`G:�Bpk0S+KVj�]�4뼽w��سU�����j���H��	������-�9D'VͷHJ�m�����A�D��M��߲��m9R lq��`7O) �4�}�3��4�>j#����
���t���x�'C�����.|��^j�g������x^��?�c�����iچ�T��~=�b=�v�)�{U�&-��U�r�R|4y�z���>�T���3��C1X%LH���� �s�؛𽎥#E̛�h�g���d�q��{�����X�M��h-C'c�uɊ�H�x�O��s{ܻ1�l����Z@�]�a�ރ���\U���&r���R��7'"<�R�m�.��	��}
����Z�ƛ�ك!��S0�߳ ��O��0i�j����Q��r	������nP���E�%y��q�-�~�$��{l��> ��;�;��H|DshC��5�U���Jg%�H�b� �w��D�&����N����{�EA&���F�K�� �{��LN��n�%�fg�V� ��D�&V�:]O�$�rF���&�/��Pݝ�6���Z(�X�L�l�8��Ҥ�<`����y�D�2V��j���(�`%$YXc&p�M= �����{���P�c}�ݮLLQ����^{JD?M�_�t��Tɪ�2W�x+}y���Xho�(�P}$�⿮W���	o-f��(�]���	'K���z�Ԝ�S1k�r�4%}Q���+e�9�� p��7)�j~%M�F�����`]\OeV
�=��Lϥ��T���I v*n�'6e��:����g��8  �FG��
�Y	;S\r7�88kَi!k���H��#�zs�GH�F��Z��ލ}���m�f�@����dU�����م�m���"o>B,Fb�@�!�w�Mv�ޟ:�U��_�]5ߘ��_;���-0�F�2M���e�_LV��px����SU���I#0��:-v;K�H��!�t�u��ǝ���6�_���H�]�K2-T"��.���U��Q[���0�	G���eث �AhkČl�׆]��/�����rt_��<��Qum�W�f�b�}�6�y��,�c��fπJ|�:vc(�sMe<�><s��u�Jl5�Փ���&�0�� w�{
wR��G���k�����E�z1/�Φ���@�> #c8w)�~v�[�r�C���
d:"���������*�</1���2��l�`����'/ ��'������Jb5݌�W��cP\��?�ٟ]��%DD��/L��#:߯�"�U>�'�C��Qp�f�L(:���jq4�Θ��yM����2����ӝ1R1럃/d��X��*��$���&�;��
P2dH���[���uGJoC��F��w?:��V�Js�Ul����<u�EiT��J�a-��ڵt�< mg�8�#�C	:����#��'�ϼ�����������\�5�u.�Ɓ���N>G5��^0�a\�s�1QDw�b���
/EFoO^w(=*��s���UQ�C���J*��R�J:P��*�:ZL>�y�_���L��>~t����u�O��~�q^�A��6
r��q(l�$9�7��UmR�1%�H�'&1�P_ɤ�B1$KY?�� �Y�1������}'��g`�� ��do�6/5Z:Y���2��s�A���Y��.�ܛ����lT��t&|�SD�L��!�6ڨV�����SW�T%a}�����E�����/��C�!]5�Φ&�g�3��5�d���l�zr�EWŤE���rΫ�FOM����$���u g�X�YS�r��d�65PoA �e�$����7�.���A���c^9�v}�XҲN��S�"�sS@1��R���K1����\ ��DG��\|Q�[�Qs�$�~9�W~�\|�J�y0�
8���"�U�8d���8�+��u��:�eǾ�0���'x��R輽5P�p�2���n��Õ� $�H_��nPXZl4�?�0��y���d�s����>9�(h�H�z�U�DԈT��H�͵��M>D9^
��A\3W��c)Րh�&����a�	>�W��D,^�4�t7�{�������i��_}W(e�¢Ut�`����m�b�*zIW�Ԯ,�BA��/��,kLѴ�����w|�N0�(��4���7������h�4�RY5�І�7�T���md^���ND��RszU�!W���g�#z��	1 �j 8m��N{�2y��O3�����"r�C&������S�!�L�a`�����L���7��+�t�*�p�-�Z�?�|Df�Q�o��փC���}�;�xP)�Rn���Ф���h3�^��z��bu��W�w�,2�C�Ļ M|�ީ#�!`���8'H����J���<E�\|ĕD���M4�Wc�/�<� �E��������&GB�-�'��
NI�n%
�#�� 
��Ru3��R��3��z㌗e�&�vp	:��ڹ�n�/V�P��Z���m�|��4
�B7S�@��j,m^���r:_�y��Y0���?���Ι�0�r��(<��(�����M%^�����BШ���Su��8�v�M(��J\�e��'�)�ֳ�Y�����~��qG�xqه���]�<Tb�Z�BF8Bɝ�mᨃh}�41;�i\2�௷����F�ϛd����<!V^��;�8d~)��$�D0���=p-5��!�:AH#�9q�~�Rez���g����s��ܦ&��d->h�ew	m
N>�|�.����5�˚�c��>%{m_�i:�\�#�e4����)S�ִ�PՄk�J���
�ҽ��\�$��sSQ>�eYt���#������q�q�'��eB:��������#�	�k�]�	��( z�H#/$�`��P�9�i�j�("��ŽR�V{�e	t���~7��]�\��E�<){l�"��A�"v68���´�k9��o1���c�\��;y�!Y��]��<v+=6�����6Y}1R���FfCH-�J���e�|�0� ��߂nS��59+�
����g����A�\�U�Շ�:�:�.�e��x8;@m��UE�R��&��5 P/���b�U�1Ymf1��%�%z4�ͪ,�4
����O9Y�,
�4i�������&j?��4*�W͊&�o�9�"�	Lv�y�GmfH���&2�{��b�9jOA���`V3��!��P��j�!�Y��0=�╋�/SI�]|	�`&]J��l����� kEmnm����We&P�H�S1�K�i�给�J���%�I�,nST��j�9��mȿ@&s��������b�5�����g/l��'�P�U��6W����>��f�?q�ǵ�Cd��t���nc�X�FO�V ��_�Z�,:�.�^Q�ǕB��E���`:�^����Ș�V��˔��	��^��F�b�QJ��X������PV^�b�����W�?db5a��a�b�f�X�z�Y�wP
2,�ܨ�����k��z�)`�v�K�#��g�q����(f�g�a��{�����>q�j�)��|�Z�+("i�V����5N�y
�����O�|��*#	���������;g�.��
���[����Q:,̊H7����f��Y|%�BY��]���#\#J�I��;��O���4���qTfh���l�s��`����X��RG�eC�?v�
Q&�Y�Z�V�H^�w'��5���L�[�K?���_��l�0��M}�y,(�m͙{�P  �/1�����+�k���0��9��Sfr�:�k&-�쬠�m$�J��|�!��f�wRi7}�gĥ�8I��Uo�'�A�$0��.����n��W;D. �/��F���A;�w��H��ͼӳ�y��{1p��i2
[��a��Y��;�3-(�x��n�Ǭ������IXuf1*�=	�$M77.�9܍��ŷe@�{������P��'�G�c��\Ƶa���N ��n�\\)�3�7��;;� ^���c�q�{�ѓ���#"�ԫ+)�ɪ3����&��6��\ �z,�U��e��>�4h�;Ȅ uXFǚ�N���@�?�Y��Z!_}u����::��L�a,R�,�s�?Ё�M�tI�߫�a��^u� �0��"���$�9������+~3) t��S��3�2KH����=\�NK�2yE L��əi���H����Ӄ^�Av-�`�Z���S�kfGS�VÓ���e�FS�yW��1Ӓ��}��j0�q�I�x��Z��9X��ڝo8�
1�=��};��	A���kp�`Q�-]���l�,��P���+@���G0���)��D�]�p�@��C/oV����R�Ĥ���6,߾N��"�Ń"�c놣x�5U|��
�٭�
�_܂>*�=�A}_��A�<�1�Y����XH^8�|��-��I��Ӂ5�Օ[g�6!��v����թ��ҒD����qaxu�"�-�H�g�a����U�J�-+/Y��S�T�)��1�-�S��1h6͕lv?��T�����Qǀ���3����b5.��6�����)���u�-4�b���t�=F8*��:��dz׈M����  W�m��m��}=�%aJ4T!���RQ�4 �[k=�%A���)@�Ņ�)�5;M��0��:}�:QTؓ��&>�p�V�>�"�Ct�]���`�]K�g?p�������8k9�����U���O#IA�%�?5�q������03�q��Ź������ڥ�n��9�{��u�9Q4:;D��7od�����rJ��	��c�M"�g�)B�l\�N]����B�.����**7ēWjO���Z�Y�u�h&��b!�흝}'�J�m��
�5��w8�����G̣�$u�+穒/�sZy��z����.�i����2Q�n(y��,S��m���hZ�=�\m���e6�p`b�{�`��Ԥ�I!�����"uL��˪e���#���
Uc�����w'���g�e���[��`���cN��C��v��M9�/ͽH־6a ;�8�wQ�{���q8I���Wlh��_	�,����ϲ%�9>� ��|,�C���g�`���B��b�Xi�QVØL�.ȧҳ�P���Vu��N"߾��x�-��0��i"fZ����d��� \D(�	��$���ޱ(jߠ���o�����0ot�����qq�I@Y\������T9�Hd֞jk��
6�L�H�by����E(�18�1[�6�K�E���䤲��\��ɲ��L�\�#Y ��/������v�)��s�ܶ:��6I���n.t�F�PPѕ��$��ӑ�(��c�5�X��f3��K������^�TV
@��B1�6W��l@��8@�[k��a0<��;x�Yt�*�=� %�\��YS�"8�^[�W��/�c�f��s^�kb��m�W{OB��a��n7�h���j���l�;���4��&!(���s�	{���f����9&ӟ��"��
c>\8���������]=�_��p��3���H�	��R����D���.0�ڿI�`����=aBl�B�P�Q��P��`�8d��Xm��ѐS=O�ƍ�1��UBf��!p�͈`��q�����tk�O�����p�Y������^R�'+mAxr��� U���m�����g(Y��^q���+��sk%";�
�l�<��ӫr�T�K��?EF�������dH��߂�eofP��s���O�qH�+�|m`஗����q(�ouɩ~G��?NI��;prkˁZ�����_��������!�C�w�t���(��/�h��U��yرI!�����<���s����-���{��#0���5N��P���gZ���Ov�Q��y69�=�I x&#<���ty�ErH8����2���O5��K�Oy3��P}x:td�$B�؞5g���!~�j�}���8����گx�I�Mc������U�Rp ���sU��!+^�:2b7�`ա�%]���~I"������b	b�'�P<�il(wh��
���.����g(��9֞�v^�+���xs�X��ML�p3���_��J2�ђAw`��|Y�UV�]�A{��<��-Mjj�ԅ:���ƺ���mlթQ��N�E����&��fq�}��2�Ta�C[)��Kb�R-��R�G���9!l`���J�W~���{wy�n ƀ�P���n�\��7Z���_�Kb�j4�V}q�R��M��.�<�T����.��F�z4�f���G��Z�n�٩�Y�~*o�Ba�l��-7�[�R�Zs�c:}d�.�K +�tlB3�*�|O`���0S�L$)����C:@��mE�m�yyʓ��9;�?�٘t閩M��h&�w>�=��B��^z�q㚨�ʬ�3��}��dp�_0�2�~xꨛn�3~7�
Q���*a�܁���h{3y<��E���:0V��� ����o�����@��uFc~�jW���R��ˆK�+�$�]�#jTqRƟ��X]i$���i��'�a�VO8��6���c�=�I���^輪&�ߋ�)_�ϱ}k�U�p�-��OO�v�w	����]Zҁ �E��Q[�i*����wQ��Q��|*�껩
��XWn?Ȇ
��0�]��W�u2�;����#:�١�ʀ�)Kq^5q0۲�t��b��k><�,�R{��῰�m�3VK�[����!��h0��`��o�����i����E��bR�E0��ig3�%:��׌�:p�%�����|$�ng���@��"?�=��*</���|]���m���I&����d`*�t��o���<�l�tN�RיG��9�{pH�뼶wzC�	�-�n�?��h��>��E0���	�9���,�[ �p 9�O(O��= 
a��}��ٯ��H�UE��r��0��<Q��V=%!2�'�U&��n�D S�.���v��GGH��;��Ԅ�=Ç��K�)��h����ڇ�&��
ת?M�3�r���=�p�P�vo�&�5@�ddБ�[�6�r��L|�kQ��ed.Į3W7�����ܓ�Vg���I���a�]��>���M����#��1��<��>��=�Ѕ�Hh� �=f���E��9D��%�"',� ����R�
�D4�<m_��Yِ�|dQXf����2	[(�\���e�����_^v�3S#���]Ey����lЕ4��v�Y���®d��a�⠺j��1LT�ɤ�S�� @���M8�Z���~����QWut���O�6]�FP���3g���&��i�)���� �5�]v/O�	e��̴�78��EC�i��`�i�V?	L٧&��	Z���!QkH�C�53ȍ�\Z���G"��=�)Q����6�����@x���%Y�1��Ѭ�6�$���f�0�J��J������\�"�0k�	�tۄ�ow�X%@��[�m�c9�S��M��߳;�uI�{��'��!`�U�X�ewz�G�*O�C�L��1މ�Wa��j��ҵz��D�2R��Pu��WI���彻*���>���~�;��vn�X5K�[��C�-c��a����"
x��`������M������X�0M"��<됺��+󎰋���X%�V�Cf�2}lū����e��]ȇ�^�?�ƬG +�v�l޹�G��sی��%hP�%�}���3��6@�p�\��	O�gDZ*ə.
@p���,Y�	��i6�c��q=��/��y�u�.4��7�A��6�#�AβRo&�?4�Q��:�s!�4�/�,�j�R$������T	C��B��z��O����h��lcJ��`Z��U�<��u�B���}4�?�d��i=3ʤ�w܌jE�Cm�!0�f���+�,i3[!?c��?=^�n�1����ŧlE1n9j�q�NN��O�k��W�=���>_�{�	����#K��m��.ˢ	K~��֣�A�o!�B�r�Q�Z� �j����3�PF;�����Ϙ�8׶�˽֟j�,���`M �ٺ���^7��V�n�1���2<|���������O�ـ۬���LhV"
�ԿH���$���8��}J�S��b��b+�JS���-��%��|u�U6'�X�]�"Fu��ӎ��@2n��z;�����#��c�hk4����Қ�Na�8]��� �a��y�(Za�x"��w�M�C�ٿ?��tS$ȭq������.PD=8�7�v���-V&¬HL9�{����zՀ�AkQN���|�����'�d��@H+�5$T-���z~Pa�s���	��DJ�/���5_�ϩ��L�7��5!5�]TЏF��$~,f=���mtE �`�%b����ym�>rx�*����r}�d��X������|AY��}�e"�%��#G��@��2Y�.݃r�R�Y5cF���M&���=��0L�m�7"v��G=�"����MK�8x�(4�HR�A�7C�����3�Z�N�ö[� R1tO4�I�+byK(�{ס0����le����A��Ц��l�2���Y����<�e5Z�-E3gC�1�Tr�=	S�F���k
В��{DSܧ+���1���D"�4XF��$�3��Q��%� �X��-T$�+Ixx��}���+&��K�@Țϒe~�'�aA��Y<;Yy0')I�����UB@�W$ۤ;���3�bk@�PN�O���R�2�y�&5���<-u.G_���vV�����k\��K,N���xQ1G�V&Ti����z.���Q
��E�0}1���W�������Q*]���ԡ̙��REv^
��$��7 ���	o�,�6�a����,��$~�gW�8��;n+0��F�Y+#�xw�b����!��N?I�	g��%b�<���8wx���Z���0�H�= �{y���#�Ը���n]K��qg�i/��r�:�ߍѾ��oc=�=�Lm(�I�_Az��Y��X㪋O��c/к�����z�,Jc̱��s�k'��E���Z�Zu���� :`7M^�O�P�K��-M�[�k"�(G4������쏷
��[���-�֤�r�x�I�U���o���ⶻhf��L���Th!m�l�]&� ����@۸$bW�sJ�qx�'a�qB���L����,`��5+otńq�{
�$�s���U1��1ls�� �h�Ù��l�y��8Ƞ��snqHB�PD� �z�S@�"��L��9�q�C�m0@��0�����٥���j����� (�iG�;/G\��׮���l��ˋ�\J䫐E��oM�muäh��7���[o����v��f��t<���r�7i�4k�
��T1�}k@���	l)��)QY̎��:�8M{,ET����V!4�]�B?:@1�Ԡ<�hw{�`s��A� ��?Gī_/����0��[� �x�	���8ac�L�}��Ф�����\:HC�aJ�d�u#	�L�8���ë�" 
�����.�c/%ߵPſ��%���Yg$�{�ťvm6�2Y���E`-m�jO�sPSCo�`�Q�S���,J��͙����˸��?�Lv�yfUЬ��_-q�۷�.�꯭E��������}9���ԇx��ⅲ�TJ�,����N��{���p�:�	jy����f2w�['�x�����^o�;-�TI��.�.�F�!�%,�j,�ӷ�x���p��Rtu���a�OEq�%W/�Un���_��ݩ���w�*��	� ˁ�4�������%�*T���5�'�,s��Q�7�8",�����G\����� 
Z�$>,2�R�2��Y,��Ϩ�æw�ˀxp�z���O
l����Ii��{��(�#�GW20��J�S|.0T d"V:�P=� Q��E��4`\Ӕ�����g��u���a�ga�a�tL�$mF��x�]�k�J�䭔�Ȭ����ۙ��]�E|z��e���d�(>�g�[��ͳ<g�9/���~�#dC��-���V����VQ���qƇ�4���AnӬ�Y�Y:�ܰ��/���)�]�*u�q��A��M�Kf,��,ui4M�%�i�΍R�c?cFf�����*,M?�P����akYhbN[��~�v�BW���d���v��Pq���N���	�Y�G`H����J���U-� ��%'	U��Q�l����yڃ�T�a�d6��!�֗�J,?-h;�	�]�h��.R��:�%:������
6���4��
`5�}H��BNه���%@��T	��nJo�+��>���X�-��2���CX�*�6�8��Cuc4�D��$�u����JE�?Sˋb���oâ�o�.��[�1m4���ߠ��2��w�W4S�pey���e�#vI�٨�O���#)���S��R!�Mڑ��UZs��R�9��f��@� T��\f�n�vZ�#�$�IX<����V���~ �V��ز
EC��d#�����6h���!C�
�H�qw���ZYV���Kz%���pPt�?+`	��lTZ��HJݛ/�A���ޗS��5�tׯ|J�JG)��}�R?�(9����1��=�v_�])��j7F��I�$t�tk��ￃ���/�>�X\�h�Lo�O#&��Z�=�fa�"��	����q��6mJPm~!�Lb���a}�v��N�f��}̋JQ#R�t#�$�d[��,~�;����`��5���c���[��n�L���s�����?�!�p�o0J��}_�[/P�O��B�s��ps�� ��+3�{�SU����7�zH2���j�g����,.�I>����6B�뀭�QM� ��F���O�xH��Gf~V��w���>Z��1+�l,5lyb	���_y���[����g��ؤ[sF���dX��|�%k�4�_��ļ���#J�SF�Z*�T�?�ec1fpƯ֧�;��SY�����k!�|��,H�F�:S�eo�Az� ��;*������@����" �&�R�k�F))z��dJ��@r����YRs*�B+�Y��a�27���`��ٔ�8Yj	�i���}f�f��Xdtf�,�����Ta����!>�����2T�AO��}�)��t�
�TUT�	�V��U,V:${�V�:8ʾZ{?�Z�י��C0��U� �C�sA�J�7␠ώ({Y�>A6��؊��������W����UK)�"�9�vƛ\����]�˂�������?�A��'p��J`/��֐K%8/���fNx�2L�n/GR������Si�y�����d����H��1�F�=�����:��D��S�x��i��+6������0�U�Z=%�醥�qA	�w�<tK:�3���iev���t�٣��i��ϋ$ԉ��v���ea2��"��a4�㬭�O����kQ�=OZǠ�4p�޺"?�p��t��'_�#I��2t-�Gދ��:)�@���'�?�[��'~A\�Vd�,
}F�3�J+��Mm�ך@V�<骹���C�bq�h�/�Gv��|�5��5k9Vqv_��\UY�����eE���c��8��x��#�1�q}յ3M�
������E�QA\���A�U��	�����(�6?��t]�*�-���+��������oE���Y�8V����"�v��L��4���@rMV[#�Bzz����~ucn���j@;���|�`'�����҃Y��䵋���'T.�H��7�1�D�i���N���nbF��_g|V�.N3�/��Bޛ�z咆���pJ؞��$�fn#^d�.���%��(g����ݢ�3�s#j���6��b�OO�e*h~�U���.����Y�R���7s��ɀڌ�]��>�؏H�e�6�X��r���;f3�6�zA�9�]�5�	�Hf:�i���R`T}LJQ��J��%����c�ﹸ�\r�l��X��K��SkS�;
�/NA+'m�]��V�(�v�I�ա{_~����b�cӝ��X���]8j�3-;,1����lO��I_-SQ��(��y� ����+Jv��1F��?��;�� ~�"���Վ������d� 2ݙfߥ���?�.�N@�"�^Q��uKy5�^$)��V|���}�h�3)��Aơ&`��OPR�D/4���~����z�Z�L�5�4��|����Eǯ����D	v�v�Y�l^�/�n��Wvza��C��g���)qz�j�t�<�����k���|'�5S g�=��1�p�ԏ(��e�aD��`��EB����znG@.����D���z�R��X���L��d@\�]'J���U�CS��;Э�2LF/��x��}��N���8N����s�չ�5��/�sn�J�J4�F�N\r��}�{zdwd�/1$�Ń�&����rcQ?�I�G0�ܿH����WzFrD��~DzD�Ⱦf�H��:~U�P��c��у�P�����R��[i7�puK��|m
<`N�z�� �85�U͜�i���N�����(?1���$oi�srt0�,�m�X��lf�rkU� ���P ;��,HGBC����:c�qs:~I����R�>��^j�T��F�5s$3ˍ�y�qn���bv����R���T�3}k��ud�b�]a�ѬF��ES����g����#֎�g#��	��E��ܼ��F^���#,��s�^�Z�^��ٶF�c�[�S6�۰8�'��^���\�*��4�Ѩ��?+�aŖ6�!,�x����1��f��?��
��|8v�xn#"��a����Ŷ�n���4��� �o:@�"�w3�f��)l��ǵ��n˗hc�@��]��X6�N�-�Mp�@ʥ�O���w�P;@�4'ix)��]��ȉ|V���L,�I��w�7����%�Y2�k�$�/�B=���¥˝�J���/����~�|�d��_>��Z/CfB�;����b�+j [=״�����w�ݼo�LJ1#Q?I�k�O�������L��؄�.�,���Z~�����4�Z�N7o3S�k�/*�;��߭F�m�2�A>�<��*��Q:�����Z3�+l�'��H����P����R���;�X����M���IU%�.�7��}���HG�M��|�l����f����ք*��ڃ�P��>Dx4K�n�F���b��V@����V���Ŀ�����F����O� 3=�s��9J!�!)v3�Y�;
�(�XBI�.�g�1��p}$>�.��tQ�u �S��i�Oe<���/xvȴpMl�8����KzK���r\G�l4]�z�5_�X�O�:�����}S��|l���YU�cٰ��n	^Y&	E�J�~�D�ԭ��:)-P�:W"3��4A7/|�ٜ�o����.�ҏ+���)�p�P�@�xA�s�q@�7\�S�]F�#2wn.,&��L���p�~J"���yz}���;�u�4{$xjز��ܓ�!�,-�R�5��A����I��H�{�B��!o�a5ՃJ��"�їgw���H��.��%eP��1�5:���s�t$�-+�~�x��e�96G맩��g)=j�]�k�q	��3�~F��W�GU���q�X9]/�������X�D�F���HZ]��Q�Sꔧ��m�M���k2D%_&���6#�R��ܫ��X!�F���w��F�+"1�K8
�L�˳��	U��$4�y����[��?�i���$R5$g�̾��
=��Zn�.�K_�UY�wY�mQ�P��WͦA�7���NA�0H̸�y�1o���Gۥ)�u?ҁ4a�� �:=����������
	0�����a=��#M�V��C˿u����M�4ax��1����]��)��#DԸ#ʓmE=Vir��%�$"y��U��)�;>r���-�E�U�l1�N𚺆����BH�����Ywk��5������d�V�G��\�K�l������V5�+[&s��t/ݕ]�tP�3,3�7,��|^bb�[�S�3�^v��_p�ھ��[�������ZU-��0׽���A��.����-�$�� 	C��Ts��!Q�U�ϳ�m#0�<��� �K&���\tU�)G�f�
U�����§�W;�����!��S��lX�����P����6Y	�%^����얖,n����q^�7�w'&Oa��f�e�8�_V� +����re�|V�B��LwX�d���)��lorWF�~
M`F���`�*���h���/�������>+hS���-��.�6����0�}��60i�A�$����7�?v&��M�iM�!D���e-�,CW��/q��n��@�y1̼�s ��ĉ���v	jS�7�~�R��JJ����,�P��|#R/��֩�b�X4�r���(����2!�0q=�j^���¸U�U��(�	�׻2��7g���i�;x���S��j�1;b^�<���z�W��])�_�QB����P��A���ID��8ۃR?2���(�0�@V~T�[Y4Io��@��}%*�BCK��#Mɼ��J�P}fŝ��'~��:A-�ۣ.�Iu~���8����:=[ߛ������=�9Q��X�N�� �q�@2h�^nMB��7.��ja�O�G*�Ax�̂�j�L>6:lhά�Ζ���©,����P)냌�,�=|@"�+)]u�l���H���=�K�i[��!_� �{�
i�0[�5�@ÕV��X��l��̻y��lv����RmU)^���,2|V���l 6}����1���7fF�q;w�s3��( ���lJ�s�b�O����������`����㨥Uuiٶ��r"� ���B>%�⺓�����!�����O]ȏh�3E�B�@�w��3�K�Y��#�qn��4fQy�����A��:�  �δ�3Ks��WJ=^�f
��hq��K8D8���D�#i?ϗ@>I��j��T@[��Aw���֝	��͏pϰ j��'H�l���pТ$�P�����s��P�p�q���
���mi�Ĉ߀}/*��f�Ӈ�?��>g|��:�͓|EB��k�,��s���3�IK�����QŽ���K#�6�*r�D�[�K/���|��
��sK�G��Q���=�	�2�_"mHKy劐�Vl�O<�k-}$��+�2i��/i4���+a�o�����\o*�_.�M�K�Lf�$wU�(-���%b��B�*zV�{I���_<���&J8,�F!� �ǰ���S��6�:�F)���9X�Y�X��|G���M�q|DXۆz^�H��Cܙ�Z�P,d���gÓtG�\%��|���bp��X�4��%�M蓩	J�'a�Di�|����֪#":��`Z�$��;q���?T��.`�+��^�:Bn���D2�����G�]0K�ځ,|�$>�������$K�RR#(P/��t� N���oM��4X�G��G�N����i;G��T��������x��5]ݪĈ����sDV����Q0.zS����`��12'y4���a� E�*���-���(�##����`�yb*SE�$�]����^*x2|��_�Mn�i�B�P�[+;�'�&����h�5	����$<���������V>�3|�&��C��tL?���O� �|+�6{�x.#�~�������y�k�-M���W��ZYF��^z�+'���3�����5~������q��j?�q�c�^n�� �/�B�QW��8��.C��'*Q�Ò��+WN��_67��T����]�k$�k0Qg9���(�C'T�S��b�a�&�3�q�,�Q��<1�L�t��xt����c�)�y�܍�=w�HJ���vM-̓��H��^�����@������DFW��g�m:J �=~o�8|�D%ݿ�Z��J-����n�ĸ��B�䠾�i4���ƌC�f�f�� |G�r�k� 㷍���3�����Ŝ*_Te��b�G�G\�6W&�鯚`�L����W�a-���S������7��V�;-I�1Uz� �Ow���E���\v��/����G\�v��ύ���u{;p������=���w_�1%H0��:&Ƴ_�]�K���B:F��	' �����5#��j�	��w�\x��]�~�"�'��mG�����
,��O�`��?
_8?�a��I!����<{�y㣀�Z��?Uy���z��MRd�?��)4�x|�*l*ǀ��dH~��ꨭK ^g�iLQ ��iW!dnj�?������h;��D��J��U�Jeˇ�"p( fp����L�+Yt��no�X�d�~�&d��]�5��
�8���+e
v{ZC|���Z�"�ߺB�:~651�/�w���3�4��*��C�S��Ğ=�a�v7`�sV'	ā����G� �ˍ5��zP��]֯a���*i=GV�����̸�,V�޼�얦�ȏ��x}�����	M�7��ש���:���v����4��<��Iޙ�����/϶(�U��=�tE��6U��>6vW�� ;h��3���SsSy��
��!���Q��&�l�iw:�7#��\��y�Z^{S�f�Y�Օ��.<�[���R��U�>s!�X�˔*�8��t\0o����d�j�RV@Ĝ�\�/^�q>f�OLq$܆W�>L	<�<A����Gc,
U=GPߙ�g�@�޷9/��u���[]ah�A	k�x���S�) �D�������Ƚ�
@��@1�'h&� ��{5��!�ݟ[/�3��	���Rڒh�K�"�V�+�q�c!H��G\���U�%�.a���֜E��������9��5�r��ãb���s`�]2|�����N��G�ɩ�:I �@�TW��T�V�`�>ox �5�n.�����V"�zLh
�.�G�	�)�M/֭V?T�I��veo�t��)<���#	l�?\u�z�:���I�*��0��!�j(/���V����و�]z������W4qn��M㤸�	��EL��^=�_!�s�UTZc3Q>��+����V"n�n�҂	Ӷ�o�W(��%sC>|�~Ϲ��x�aRD��Z���o�p�$��sG�:c�tKc ��R;���H��뫴�����	�/��6g�V/���0[;Fq�a��P;`Z�V�nE�J�gp���ԓ�z��ڒ�����a@��Q��� �YglKd7�2�]��Il��c��{�7�P������C�b��"��k�����ޤ<#�ʴ����騉k�D�$�nu�?ɒI��p6H�A^y�:^���(gjdg��I��	]7�C����e�ԃ�E"3d.5H�ӕd^ JWF �����nY��eC۾��̱])��2�t5�:{��������ɋ
�����k;Mg�)��3�$�N��	Kx���[�$��wEy��%��X�J�����Sz��^�mh M_f�vV�����I"��D0�C�L��az� �+><]:��v�8Y���@��6��[����>��d�J��g�$�|�wpO���Sk>�t�78Ӛ~f��3s�K��/-*���w�ޠ
 aq{P�\dۿ���{ڏ���|5��AA}��1D��� �oM��-�4bWr%I���KF�Epb9섃i�����Q�'�A3�y$ZbI�t���#�н=��s%v:��3��j;&[>�Na6+�$�1��GP���@�� ����H�YӀ[`�a)��B�N7����6���Z���k�$�!j'9�L)�(�u����؀�o��	�mUcsae�O�ô@lAM���!��}\��/����x����	$Hhu[W���¬q͐�$6,�9�Ëά=�U�bJGl�(�!��� cL���0mX���?�̶	��	ѭ��c/[��˹U#.( ��|�2Pf(.;�u���s>��I�z��$�ɇb$v��y��=�ַ6������?y��$ـQ���y�t4;��Nf$���,�~����������͹46S��Lf6��r>��;����&6o����p^��%5�Pg�v^�����e�O�/�p��K�|��T]청���Գ�6��$�eD�E���]��G��I_�B{�En��QJ�z�lP��qOJ���ڈ.��Ղ�m���I�m@�``��.2g{y�f�T�V �,��M�J?V?�E�Qn�M�������/�g:��rpJ\M�lHqm�n��jZ@1����+
���P2�/���>'j��+�����DK�Jx�O����"��j�xПЕk@;����u�6�{ @CJ�d�-ZC٣�YF@y�0�����\��c6��VO�������I��X�2��������z��R���z͏#|��,�t�}�������b��dL�i��y2�T�3�	�6a��^�,D}K��ޔ��/���n�fw��x��P��VQ�厛A0]�]δ锶�_�	o� D��������o�Y_�I���[�c��a���J>��� ����*#�=���%��-l\dY@>��DF2�?ۅ��.�J��j�K|<�����)����\���.��kU��ɩerG���x����J�n�bx=v��X��\�i<�3��M`7_����=]c���XF�*ӷ� 屉�y�*:U~�B���*����|����ZP���?�+��l;���y�6tK̦�u_/Z��sl���T���>��Jj�	@\�w��&�����2{K���(�~�w�-�ű9����K�U[6�����K(��3��a���q*�@���>d>z�����gK��E��>j7o�A����lB�x�x�\�����l�h�������9ҩ��s�����(Y���9eKu��9�8�H�h�������8�j1`�Ɂ���e��'�����̰��ZB8Bk�|?Q�(�{3ѷ̐���<�M|n��l21�Ǎ+7�����M�>��-�?a���^|����)3���y��|C~V�E�YE����#ڊrz6x��5�E�I��j:X�n�3kL����y����>\�%��� ����z�������eB{�D�X_�5K�q�s����\ѭ�'ϊ"����,�F���|D�K`���@��.���!Μ֭�/��~� �x�V���Y�:Ej_�"�����,�?�.�U��nϪ����#�8;�h�!xџK�����y�:z��t��L/fIҿ�8˄S7sDbϸq�2����l(�A|vy�؉�$+��U�o��ޓ��[0��"�[i$ϖO�	N���:`8N��R�޵��,Ulp��d=��n�����.�]U&��9�%��TM�
��W�0D�r�c�����^�l��Ye�K�AUy�u$����6�&�YFV�x�֐숸2�L=����eb��:��х�T�5��/��PRV+%�@���)�_�L,��v�-Y�20�������v��;�|ǿ�o��W���I3�[P�N�F��;�0F==Ɏd�"�+��<�a�dT�{�E����*�:Dw�Е+oIw�����13���ug��"��c�#
/���K`�G������X��'>���#si�Ζ�I�u��q������NZJ���,�&h��o"Ǳp���H�4{�XX�Þ�6
G�̝�Ej�W�N�P�� ������Ɨ�����JA��Τ�� �D����7��D�~ɤsG������&.\Eh�[�?�q0��/�#����D=(�f�j�ߨ3��!�^a��/���lf ��C)_�ԍow8��B�e�ɦ~^K��7f�'2����J���9O�'1��z��=>Zۉ�<�i�G��<�#�Y�V�d[���a���T)�3=��J�<7���f�;2���U�x�����)]4�f-ȭu�	��RI�:i�W6v���n�~��`�����o�i���9\���-
WA6�K_��]�|�(o�َ %�gv;a;94`��)�]D0�*�7���z!��}O�b5�~S�3����2=��Vqmށ���.K_<��~V��
�a��/�!�*¯t1��cf���ǒU��#�!���|�`�g�w�{��{�q!�B�����p����b�P�`}mf���,jR��J��Q$��3�4O�C*�̇8<�)�?rȪ�^�Z�@c�Q�3Or��[C��1�Ё�I��E��'�r8����zz@�dSbM`���t���{��B�N�2�z�)`1�	C��Iœ�H�XIL��>�����|�M֋�E-��?�^��y��h$%��w�!͔�Ϙ�L�#��p��B�����d��c'BȑRȎ���,��f��U+k�@_t��_�RN�� �YiF��L'�ΫR��ȿ�)�#���yC0��ˮvZ
�L-���vgZ�;�'�/J%n��Yz�H0���ܿ��z�0=Y$�p|��4��W&���ֽ�v�[)��8��!Z��]_��5�� ��:��%Vh�sp��%�H�N&D��LY���� ��i(���"먙�q����JS����3�H��R�jo����:6��R}�tɊ�0�G�X���y�>p�b}��z���ק�/ڶ�g	�|G$�v���ɍ�Ĳ?����<y/n�x�g1�(91��V5D�L��Nt��MWRp 3QF�m}|^yͅ�cz�0-w�}����9�V�P�I;��F��+NzT�Ӂl_U3�n��Ra�Ϫ~fʠ��ȅ��Uw�������vb�A0O,�S���Ū5LW������>��Z$-�ڷ������;K���<�F7��ה���g�qܕ,wJƓ!�Q���> @�"�s��׉-I��.:�?�@��!���a��U%� T}��z8 "�9)S���?p���B��=�A��j?6�-��"�8)1+�Q��Nӊ���C>��B��q�+<��(�IjUZ���>]�lLU�;�!����7wiG��2�$SuN��!�y���k����Fj��z�p��ö�������Q���G��7b���n���h�l�.1NVm�L�͗u�c8U��B���[&�5�S�qʼ�=���)�FP�Mc�#�б���4���_wދ��+���	�c���.�m��~7�/5�rZ���q����fn�h��#��q��a�W�ɒ�iK��@�#�|�'{������k&e.�U$:�'am� �������3A.�����M7�ѫ��&&Qf!9�yN� �}Ǽ��{�1"���0\�{�Y�Q�0U[7��<
D�\'gc�(t�ՠ��O*|���{9l�E��D�qi��i��_�~���w�
��%�	���A�W��� &��y�D�����:�����1�, f\ʀ�&|�ǽ���c���
�"R�a;B��+��N���x&�DG�~�'Vb�u΃e���݆��(��*�������h�\*G/�i�Z� e�L/�VP�m&*.è�#���hM��/�Ì�p�'A�����%���<���gb��)��[,�L���[c,�Nu�8��E�t��yV��)�n���$٩.�"���m���2~]���()}&E-`���G%����8 :h�~�=�`�TA��Q8e��=�͚��d���m��P��o)�g�6b��`M�Ѯ���(EfC�+��8"'�[M���b���Y���ٰ>@?�_Sp>��M*�f�{�6;خ�-S(��p�i��:�p��}���I�<G��I��Y=\��2����lX\�rO�]�� /�l	��|(o�첼�&��~2I�e�%��>�h����X?�ݰ���G�|kd�t�k����_���ժ��rL���5�Z�_rE�NόՊi��cb0c~�h��hH <d��*sUH��Ɇ�'�n�d��=�R|׺T�q/�=N�f9M�^��^W��(!�����t�E�������<�b�M�p=8��4n����B���/����s�%I(��	R)`�P�6�L._�e�鞎��?}yr��]k6#.
���M��w)�3%k�1$o^60�y���L���e�})y�����ţ
nD��K|�������R��"�ь���6D���7��4,��s��|�G�U$�hvlv�\]'���)d@퀚MT P �}Ѕ�OGj�j���o[rj��C�|E�k4�9�AD���f�i�gj��~�k�`	GAt�1���,[���{�'��n���p�uk%w|Z������OmL�m�+�#�#Q�T�P�`��5�����i�Ҧ:������$�;K�1�{�Ĺѓ�G���W���?����5�Z�IAZKn'%K�	,^�W�o�-W=Z�	j�\F1�UY�(H��5LX�'��~iU*����Y�$ۣ�w1�@z��c�L&.��f��.ھ5|�X.�?0�z���d�_���=� [�r7h�\��Ue�QYB��F�aK�r�Q�at�/�%B&�N���k7�w1ּ=Ml$�&�j3� ��7g��q�)"^��ӓ�������V5dt��ig��/��h:����FA&v�&������z�qGG��n�n�<�$ڞ������٦�=}�Ev��FJ������j�*�ށ���9\)�h�yL$���F� ��s�M��s�薒?�	.��N\����3��n�}��w��T?s�W��Nȶ���P�[Aߵ��PD|��|�M;��CY/�u\n��2����9��d�U�V��J����D�C/�]�ׅ8�ℷ���G7t<b|b�����2�əA��B�Ź�D��Z���f��څ�������l��w�f��L�y!$��J"Jⵑ���8�k��ۼ���N���C�f��}���h�|\KBaͅ`��}!����*�d��J�/�E�e�ĪC��i�}|���OB����79ܢ���#]��2T���	�c����{/�A/o��<0�d�^xkg3��~9k�\/��G.�+V�("U�����M��W:B�f�@J�m����d��F+GB��oIh4��s������n;��H� R�j�=���º%��T�^�{�Υ�/âmM>�����Gl�G��Pl��W_�# ��V�<�X�E�����]\���y�o��ۚr_��5j���_�)+<~�kI@`_a��a��b��|Ra��lxs��s�p�a�ևN])��?� ��(������6}�;��x$@q�y���&q~���r�%sA��S���G��
J?؃�R��bJIԭ�r��W�ѡ죖�������N���f;BC�۵!C�I��{���7	�7`���j�G�~0��\9��u�f�����8��~v���M�ȉ����P�?"�BW��ɍ�	�`���5�n�d5�V`�T3+���4���|_�L�z���7K{��3�9,{��C���̾���X�2���[7ʅl��@ɔ�� J�z�!a���H��O�}$E�k���%k ����I��CK�TR �[�D.��x�@�Ʉİ.쥼�vp�y�Q�a��$���<�8=yK�۰�g\y�`ap�H��:�1$�ߧ�U�*��6�+�����C�)/7�������4�Zl̮��+�*��Wy���+ :A�-H�Q�>NV�U�x�s`�-B�+�ܑ& �n�A�=�:S>��d�97��Xt2i7�����Q	�5��w���\�!��kV�z��6Ր�$����%U�@�&������,LC)QҭH�:a5NHག�ֹ�vKI>�a4��i(uf��ן�|��Wl��t��v$tĆ�_䆖���V�fbr}�ڦ-�pO������q����߀oX��W����)�����Y� OTh�/�����֟?�߀X&�78��^kb��:�����Qq�G<�N���A.>�Iɕ�r��c|�y�iM��2�Dm�Q��s9�̆oW��*���זn]ν�(��(�h�+Y-I260-B�T�-�<ac/6#JIe����	�K$i�s	�-6I�r��u�YF	I������.#��Vm �c:ԠӞ���'�@"�߀��U���e���bbL�n��}iC[���"'�X�ͨ���'���1O�;�_D��)��rF`���u��5��� �I5���\ P~wڔXԎ�1;�@�Ji[�W0;���e�=/��X�s�D�I���Ʃ�����4ν�B2w�������[Ժ~�
X2!���X�E=��~�2���"4�U4.p�0Y/�>O�0%�{���]Î��c�m�����2k�V���WG-�����Ez��$O�A^����g<�Պ2Л籢��4f[�u��i.��@`܃Q�.�:�HI�5��|���Z�����?
4������)�"8��sq�p�̈`CG��޲��^��A���u����P��Dvb[���T�f��Qe���7V�lh�@��X"���Q�bU��&+S�$��N����*X	L9���I��NQ�y�GI�c`�k|��kF�X>�+V�:6�����A���*���;�˿�EX[Bj?�����ӌ�Q�b�e�>�y8�r�H�+{jٛ绖����_��s�H�$�2��t�,�-�ʅՃk��"yTg7@I��]�������O�r� K{�?�2`2.w���7�|���t2v �J�mG�0)��,K������+��k�������ܒ��67��,h��+���ug;!��'gµ9���qh'�s��H���?.3�q��*�G��a�=����e�mM]�1$�Mų BN_���r�=��}R��'�枘K� � No�ӽ���;S��q8���J�ӡG�Mz;q*i(@ 6N�.+X�������s��:ǢG�����^]
�O��美��v{E{q��Puw���n�T���}���L���_�u�����y
��d	|�z�y-u��m�� Ԭc�M�fjԤ��n8Y�����,��fX��R}�0}�ǩKҮ������d��c�~FC��W��^Wf�!_�VӅ?�-tF^K�z�����]kY7��5F�����`�jW}�X��0��Qc��T�!9J�-*h�����,�j]wH� c,E�i`WȉB 1���V�p���4��瘭"Ey��N�̔iUAۛ����b%ׄrw��(�ȳk�(���o]�eF��{�H_p�S�dK��B���/�-`�"���n���HD��9�
�ɼ�^0 ��X� ��PYԩs�����TOT�K��}�=��/.5l��d�',�8�e�����`=�C�k�)nL�H{ꖻ�T����N$�}(i�*At0�Iog��bn���v���1Q|�XE�½��:���Q��e<;�0��D�JC�,�����q����5����m�B~�SO��!��p�E=]���a���f^@R��ïKv,
���3�3��2���/zR˃Y�0YZQ7��}���ް����|�v /�(;=D�4��}�2����n��vW&'���FT?Ȍ�h��:\�h5�� ���q���J �	��BJ>��la��	�~M3T��:4���a&����fY����0_&]�0`�k|}=vZx$�G�L��P%,�}V�:XW5�1e�Z��兽Kf3���!zmE3#_�ӡh��ç'�ղ�� g�̇օ�g�]� -P�̫��0%o�'���Q��?��Bf&o/#�WV�m���0�W0�qr3���~�f�g�t�pΕ�XW@�9c�Hnɞ4pzɮ��gz�����MɶX���w�		C;F������6����{�aFU��gٓ��|J7M�a؋A؄�sꯣj?�?E��o��p�S	���L���������_=Ȃ�v�˛���*B�0��e�o��]�N�\X�lv���*@��iw���ϧ�BO��I���gY,|-���8�Q��.좪4D��M&
<�f�֟���a��`�wG����e,�^�P,��47[������L��A��v��ʭ��޻s,O=��Ua��8KZ�BXf�+�i�N� A ]����P�Rq&{�"<9]�*�+��}e���� ��?2�4�1C�h������ˡ�L{�c���������CAq��#O��G�A3�[��)��z_�Ż��g�$��9����S��D,�z�pӒB�(H3lox�J�.>}�\�=�O�[Raz���!q�:P��nj�[;	���J؟�^���e1��}Vv����CI��d>
�*C��%BzF�Ɣ#�>{/DS���l���d�j+Jyc'i��񚧀c?�E�ד��*�c�yav6�h�E�s9�e#d������~�"+�[\�4��Ap�6T�G�%�*����7�u�,�ٰOdC?�^��̊�G���V�hdP?�7� ���I�~`�kP����W���x�K�jm+��^\��Q9:;�x��Q�0�W�F�)���e����[�hӚ�1@�)Ee~Hbh���)�����}F�[%>U
�Q���;_�π�ߦ3r���ɦ�~U;��=)�S�\[s�G�l�-hH��&�M�(+o�oG7�%�}ίC�4XN8 ����Gu�+щ��׋[��Zu?ё����ְC���4���u��תa�e�!f��*��Qc�� ���������U���ᒿ����ԇ��\������I/�N[�E�{�	��=mӝDS��r8�sY�p���#<|�ﲜJ�]�&��Y�+��%[�FX^~�Ͽ4f��r�!~+L|v qf��('�G���h۟n�o�S���Ƽ���Ҩ�����1n-��`3 ���ԭ*�hOe|�{D��N��E��W0���-���Pd��t�2@�A׀a�-�z�ҧ�W���OG?���쎓���uוy��Lє�Ԭ�2�|-M^S�~��;�/1R	���z���+>zFi��`���&�@��s<@���2��B�y0��j+����g5��%�+�h���z���7��З9e���0Æ������\�+��jn�xX.5A�j�H�]}�y;��W�Bb�T�K��͐�-�ih���
B���%|�}P��1X95Q����~qA��8�Z;�O
��l�g��x���׮���?bY�C��F�3}��t�S�Oj*MY�ǀ��n����ғ?"vi$��珻�? C���h���09:ʊڲ����&�̼������G�(����"���B�*Z W=L����e|���>��A��{���E y����$�C���P�ЍL1R��1rE�n��K޵<{d+^�L�LAg���p��	B�z��#��y�?� �2��FA�he7<�u���g��w��r�����kq�B��J���";%d��X��|�C�dƟ����'�����u�3���@��g�A/��gԡ0�ww乱}�0�r���*��\���
��@���k=pE�e4��.�Q�p�j�c%-�x�����Ĩ��;���Ź05z7�I�Μ�=q�����x�,�;S�B������:mj�l`x�v��t5f��S�I�t������K�\�����wq�M���ɟg�?_�4�G?r��'�7N�KE��G�&2/��@�uoe�a68��ſՎ!PX{KzWPR�Y�:��]�����(�[��}��7&ad +{0�S-��#����v��v�W(fɰ�L�4xl
���?��`��VJ���Y:��V��?��o5_!9��D���g��H�=�S�N�c� X�X~HU�ˇ�>�-��?11֘L��gu�
���kQ� ����)�[D���5<�pu��15��X�F�L_����M:zi|��d�AG9$y� ����k���{<5wTh^�b�����v=��4B�����8�b�o���v��Cx�/K�Y�#5�Z�䩪$���R��`D��Ox���m�n��`��\���G�{|�	�4[ц�pwHݵ횀�[+��&
�D�����h������J</��k���/���*�6��؞���@��+��٧�ho^��d�O4+�
I�}~B+��h���H��=4�Z,Z���Y��B�op�J�e�����V+Ǌ��C�YfuX���s: �F@��齯�W{Yp�ID�vhof�Cc�q�E�)��I�@�F��b]�':��LȦ�]-��P��n�Z/x�r�b)Yh��ÔMd�N!�rs
�wV
{�����W�y\"]"ʕUZC��\N��n�gĵ9��8]��jgc�Y!@��u������9ݧ{^��B�'g0\LY�����g\�'��c�O0�u�@|��(� �Ĳ��i/�d!�cО���7��{�bÒMtO�| �� �Mi`L��$�Dd3o�JE)��bs��l����mV�$`)�k��ݜ@ƖXXA���ϷOx�iJ3M���Q	K['U_�q���/F����8k�j�j����I~܋钙M�����7��;П9r��F/X׆�s1�
_X������R��դ��%@���1���g��rN�A|sO�W�+�V��{U.�<��=��p���
��޵�}�z:��Z��1�:�R8aj@�;>�Y���\��	P6K��6��;�'�gJ�+G5'�� �@6d�A��J�peИh"��K�tΆW���<��Z�w�/.7P�4f��t#�?�g�������M�qI�G�BP��_cP���9%G'L����i3�b8�j\��u���5�
���`:�,�)�L�{D�b�a,Y�4�Fv�]�9����ā��(C$�/�d�|I��|�V�ꕰt��eҔ���X~*);�DU�wz�B+�T�\7��Xh��F�C���"ΰ�c�X��يj]������?���O6�[�/����\���]��@���9�'��dQ�*a($��:����t�.42^%{���[�-�[�6O�������F�6kY�t��	��@�m��J2�vq���/	S�x�o��.`��|jF,6�K��R�.������}�����ʹ;���K����?�e��n���[��r�Z�6En���Q=~�r+�7�6�`���_{�^u.GB���X[�dO�X���H��v�dt=�Tl�4JC�wف�����`�T�P�
����/Uܢ�>���M���
ҋ�(�!��߫�)��S�h�16���l�P�q4�y�������`:ْ�L^c�@9V��j�%�?�Z ����N��S�Z�ϭ�6�oIb��b�-�n�<�W�G��1�i��+i;�r�Y���l����`r���ϝ�*�YV�W/L���G,�]������Q�W��!�h3_�R�;��2O9/�ϸ�C7���+L)(c��Z���6���s ��Q�� ƨx���׶�>\�1A�WFa�\�I>��xY����-kib,��Q$x/���n?@*aM��u�"�[����W�(R9���AL�ݬ^��Ĺ�'���ƌ���boC@�q��&n!\m�Zk�se�E������g��	�Lي�a��g&�඾��+/����:-685ZMFBFM,Eq���I������ ���1��z��X0v�EG�9��اn��T{ȱ��D�I�} m�]�*�5X#?W7�I@��M_f�<�l_�$���Gf��y߾v�k�dtݨD��%
�ք:َ���8o,�ΫyjF�UВ;e�-�{c��0�9yx7�Ⱦ��9���'���� 9:fD�D=֔��ga�Y��â6�y�4��t#�9F1��T衽 R}.�8�1��sw�����?-��(z}�����sM>��g30��T��� ״&܄��N݂���W\���xyD�Y^�8�B������eX��5r���i�J��9��L`;s��н��0� >C�	��k/^ gB���Z@�Sd�>����`��qGW[&\jٰ�s�6��9 ��e�҅{4Td��5$���9�����ĥ'�BWϚ��QF�L?��7���tJ���	ꜷ��3i��[Ҙ���ub)��m�z��˓�.b�lh|���� c�J���&m�v͏����0�G�^]��#�䠝1���k��=4g��q�E޼;]�	��CՏPA�������}���	�:wI��xHO�Zœ�
���r�
�F�L|�-*Fx�S}���a�e��ݼƢt0��kB�>_����ҙ��j{���o���W�&ʐԖ,q!�dcoL&k��1ҁ]��f��wJ�,@h�'p_	D�ɓ�?��O���7J��+�"=�wfDp�n�u�6��;-<�3ˏ�2rk)�,�
��ε� ~�x��3����E0�^R�h��n!��}{��WA�q�~Q���k(��4Y+�5$��-
��ba��F������"mMA�>�MHH��b��S��_��	hU�|a,.���vX �+o��<y���pS�r����T�.F��LA��;�<Q�@���XnJV����.7�#l�	C��h�ܷ��m���n(�7Zƍ�xصp��Nˎ��ݑT���� ϊ�[#��MItc�ǘH�4;ǁUWy��T̠���V�9��Z��~�k@ކd���J�Gu�M�.�)}�Y�4�s�3�}���W#]��"Ξ?�9[��DL�Eó����~�q)U�<ڀ��M�{����,VƋ,}{�-��ٳs�a����[������(U?��
%����wq95
*��a���U�р�ovŧF���2$e����`�A�8W�%<o�}��y<��H������6��x�n��_��r����Zdq(�h���D��"3
ǥ EQ����������}���R�}�WCo�Q���D.�"jQ�^t1N>�����k�����b6$��_K�rR�v����P��J�d���"�i��5=�a����n���=I���S)u|l;��~�B�Cc򃄀����ڈ�2n:ȲB�F$a���#��}q����Ff�&������L>
b���#u�wڟ��x1eY��ObȌ
��f�Ч'K���ؿb:��z�pͻ���0	�K6@ ���i=W�1��a?s�)<@G\2.�w��Ľ���a�`yUE��S���QN\(�0s���L��]8B=�l�K�����y�r��F�Q�q�p�Ixw���Q�����~��KЌ<xN���2�����(G+�3i� ��f�)�D𥉉F@�z�0�?��5��d��@� zѡ�J�{/����R%�"���F�a��X�����0��@�0aZ�A@���
�>�� �'DR7�V�@8��D�E�Gi1�8�ɁZ6�3�/qoWtg��#�Fe�R��
J)����5�;"�{ΝF_���!G?�NR2�1*bc��^"%C:6�'���w�^�r��I�{fS�-���2�Ƿ�l74�Mߏߒ��A��%<	�'Vp��ڗl�7��W��Q���v��
�/�Xk�3����6��`���\+X=J�^`�8�1wR��x� �����"1s�����ʛgQ�)nt��V]���p|�8s���Yxi���b�N�5
��<�����N����;��nu��>θuZNY'eǚ����U�:
6 m�㬙�Њ�)H�,�����Ffv.FM�8��<�w�J�5RJ���-�ύ���쬾;rI���7"�|��u:dr�i�W��b}�ˤ�W�:@�2�y~c���:�b�����C�T������Q�;E���ST>�qI���ӆ�Ly+/P��j0Y�*	iM�.r��9�}��:6������p�\�Auo��{��cH� ޒ_��5~��֍�k3����Fߦ 㵊�z�F�|v�:ctW���
C^��o0�|���1s�]�/9i��x���[DpBgj�&vb�V��FZ��	B�lQ�������P�˨=�f�*������5R���.����K�(>�P�Ru�F�u܎t{�,�M7�x5����Ųn�S�0�D�t�.�B>�v��#��bt(K��,!�éJҿ+Uaڹ=k ���=GHH���D��W݅����m�՜6cX���X-ݩ8��D����I�T�=&���O?���OrB�/�ã��/^��e3�oI6���ӳ��6����8� ��>�B�[�դ���ĦwE��_׿�O��j�7��<��Xޥ��ľ$�sT�&-����H���UT�l����Y�ٰN�BR�¬�7
Fq���LV�u��4L$G5Y}	F�ȭ3,�'�V$Sn�B}A�� �_��$^���K�����/'�����,�$�`a׷⬲6��h���2Kq.G��s�>����*��I�ċ�`��N��Q��0�,��HH���������.�B�$�O�/�?���OR�������=!������t�Nl�՗�>�����@��a��k��������<�;�ʾ�yǨ��o�J)�2G���ȏu��.�P�[��*>1m�d�2�Sv/>�vb��q �����?i�����:OQ�o� ;�N;j9&�-�08^�1@I��U^	�E9����V�OM\R���Q���#�84F�k
g��I����`~��`ʰآWŻ9���P� 1��U_{M-��;o����A��C�~}u�.=�&�)��#��������U"���*�U%2�	CYط���q��'����W��5�d�'�]��BH����״E�]6!�89��`�
�%���x��m���~�Kא;�zyzqx]�;�(�ace\�I)��4۱ $�ON���G���UUI�{NX#��[%ڛ~<}1�����Xe�SH�y�+5N p�OU��.�4R�U��� �������qfty�?н�Q:�C&�KO�H4�祋r�>���:�*T�4��bk?����Y3M�HR�R���\�[��ל��o��ʈy�� ȫ2Z��h�?�����0��
'X�i{�6�&����!�����&fǋS�-R^��Y�ꈐ+���]�����,�
�J%�G������m��8����NI�]JL7D��7�8�'����1Y�s����׼��ʆэG�^���$�z� "D���^=���nV�FG���K���!�9�/⭟hn8��B�C�GP'�;�c۸݇���:�'�_�/�+YB�oh���BXcV�������m$\Ex�n��Y���E@������;��T��@,+��`%��z2i,�R�Y�#��t5tƐ)��S2�_k������j��.4��t�{|�,���&�n��Z�H��p��=��ˢ¸Z�i�5r�}�B��j����U>Y��s"�{�� �4P|��g�AB�J�0!H�e��j����S����-�"Y�������g�ޥ)��&�#��حPM7-M�0�T�@0�a����VF����B��Hũ�i��=.s�?}n}�傑��u���}��?�ꤦ���!��lUs,���W?J�$��tw��^Gd�\��Q�1Z�0�LoS�/���3�a<m���c��:�Y��:�P�y���p�3�P��&�5�LG�.�3��h��5�=u��G�~v��k��U��B.���G@n9ţFw��9�?�2���@���+��z�*e�j������\琉�6�x��S�v��`M��-ڂ��7]�q7(�`��[*��\��@A#y�w!�{���0�'�_����Bq؁�g(3&[_��
"�Zՙ2�:�
�]��]��oBj!В�N��l����;Ռ�#��	k\�{�<�(ڽ����pރ��.��8����U8|��4	1�<�Y'�yC9��ե �ً$��y�Y'�w��v�ӾD�Ē�Gzʹ��%)=6/���jʝ*|u����0�R'�ʶ��1���oŌ������ϞD��A,�����_e���z�N)YK�DC�j!w�b���wA��T�1�9L�l��-�2K���6�Ͷ��=:�6r=D��XܰӬJ�5�沂.�*���Le�T�am=��ȯ �iO�:�Ϳ��S�B��JN�/�,�v��6r����tΥï�ʃH��"[7���g���?'a��D��k�@����fz�x��ZG���k�n�1�-鷾l����N�A�@|عX���4���|�` J�w$�Z�4�>�X�u�s^��A���'�l�c���m:f��1T�W�Ae!�-�X2榸�G�+��7�����[XZ5����N��D@�E�i�:x� 9](��Y�CY�^��ヺ�Z��& _��<�����::��\�2��h�2�:��c�$ߞ�����l��=E$�� j�w4��o��|��^��+W��2N�i��`L��҅~��=t�NyɄ��0}`o����m|�0�X��ļv�`A)�䞟�r��Dl�(fA�U�r�^�s���֠A���}�Kd�3�;#=�RB�펕\��k�5,ŀ���6*ql3�8������~z8?�h��*�O��`+�I��*���o!�&~j��Y��x���G��}*O�=�-⯏��G�� �*��#�4��z'"{���"��η6V�h ��_��2�;o�c�l��
2B��c��Z�/$��`vsƘg6$:�-��S������+�h9�x+�k�_�����jS��J5g(\�����)�H&��&k����'���.��$�u�o�J�����ߩq�~6?��|��g�o��dQ�����,QR|I���g=�U�6� �xU�S���P�c�o<��c(Y���m DX~뷼�B�ze�-p?�����C7|+��"($��aH�u����\=O��������yܽ�u��_�6D�o�$�Φ#G4bϓk�,[�|ET8?GUM������2L��C�R����jϖ�*�`�N�"Rǒj*��TΘ4+�^b+5�V$=n����o|��OѬ/b/�A��Y��%�'� ��2���}C�5��9�w�� �/�����!�W0�����h~'M�����	Cy�V�r�;�ڌ�=����M冶�?���q�V��s����4.姖7�>^��K׊8�]�ޠ�����@�f�g
,sE焆��I7t���s��9�'�s�[ܯ���.:�'J<NaRۓIx��
0�w�N�x���AP���Or,��j�'�1.m���x�
!���ro@7�L�Iy�r(p��vv��� �_`�E����{���� �;+�;xj�ڟ�xct�f��;Ie!|׌�:�H��.uMR�����i�m�n)�oƏM3엚�Y1-L��(��)$=�t.�kd�_|�l(iW�u��IC����s��,CWo�h$&���S���C|�!|m�xS��:!�184���Ѷ��R�p����L�U~�R��J�<ёzX��l���5�{%j	a}���t"��Y�Z��N��W0�7�_"��6U�(�^����\�nB����y@��T֧#}_q��������~��'�w4�˕�`I�� �CϽK��n���w0l@8����,�v�-A����FzOK�����5���R�oy��%�Z��qO5�j�LV�~�;8��Z��?v
z���M�����-B���y��%�0`�Տ�C(��Va����A�����שlZ4��I��{O���)��⶝�Κ8��1�]��E�=5;H~����۸��N�o��F����y�F����(�K:�B���L�[ ,�dnn��D3��2G7B����t��>Pq%�3˻H5�æZR������ �;��\%�V+l�|a�#����d�J�铁RFàv���8�� �����N����<`C��J�s�~��l�֯
�X2֑�0��Y�y�<Λ����LI�t�!e�/�������퓙3ߞ
36�#��<W�k�a9�o�wsLj�`3�2�n:��gؠ��zW">�ơg%#(������ �@T�d�:�������@8'�)<�!�{���Sg�D���w=�{ԘYU^Q����Ѱ,�w&�t?j:���E���Y����4n'�v����#����6�ɜ�)щ��	D�^�cv.0�ߩ�W�����':�l��X��9�K�^G��@���,��L3]�[R��7SW٦\f�$����6���N��NWc�n��\�4�,mJJ[�ͨ��|��Dh����c���Qj�����f���$=�pdd�;�n�*��{��d=��P>zX
�!�e���#P{K� ����d+��fEP� ޚe��ϪP��S�p�ja"�PÆH�1�(����MԞ��Xj��~��ۇ���σ���r��<.��2r·�����d�R�T�.P�������֋�,�r���A�y��R�r�G�8v���(�H�� �}����Yfi��2럔��r{ee �y??�ސz�P}�H���'�O����;b��'�2n��Y��J`V�͹V$��mў�R�*Mph�h�_�U��~c�o�~*��@U���f����t���fM����h��wv�9� n�+��1����[��o �ZER[���1~��"�����U���R�k_Q��m�?S���sKs�������tQv�����rO�m�Εxݥ�$v�~��������aX�5c���5�:.� ���.��c^�n��g��������gjQ.�^�	k�iQȦࣚ+�p�hLꄍifa������#+٤%IP_F���C���+�Am
��P��%��� �|vd�L|���0��y�)E.��u}+�m��'-���w#����a�.�nv��w�]����"YɁ1�����"�qh���O��3Ekc�u��Ặc�k��"UM��!� S,�d�}L}�*F����rR!�t�X=��Uꅿ�ε۪�.y�uIS��UA���(&?[��DW�<��M��XT��@���/2��_O��#j�Oq	~,�r��C��]B���a]u�*��#@�ҋ����n�d�^p<��!2�d�����i�b��B����_�4�i=*ƽ&{RP�.b�#�33W�FRC���M�P��z���nk�>����	Y���ɸ)\ �a�,���x<r�Z�Հ���oV��<MI^*�js#h���۴�" �rSE�DP����"[���ޒȀ��}�]4����ֱ*��hN\��+�m��4G�k���Z��,T6%�7��6�[H�Ԓ�cQ<�ƷFn���6�
��<���1�el̂r#�Ѩ���Gb��	l�� LX�Z}6B���;�+�,F��LA��?���\P�8���BI��djx6|�/�Ŵr6�H��ps�'��=N��-%���t�yI�dU��կ�������7pWm��g����Bi��-�5Rt���g�C3���b�����(DY���%��4���X
T`t��+�p�S�@�
����(Y�C�G%�\�W7�9?xt٘�L*��)��,�g�y{�4�Ky�xf�?H� G���K@Ajn�~,M�袸&������u����^K��Ff�s!�w��0���-��6�~��\~�<~x�{T�Z����c���������s�����H��L��Cd��<���'m[������t��PaE�SӢ����3o4F�Ó�[�{�l�09L����X�jm+Ố�S?����5���M��m�]��3�/cᖣ�Ɋ��.�0�NI�Q�X�z��'�>�{<�5���k
[�/L�X�BJ�m�P��[�L��,vR�q�+�Iy�����>��59�6�[��ӕ��&s��?�-xiz6�+����a�{Gt�{.1$�j=������Me��S�@�[C|4MC�a��假���Uv[8 Ɏ\�R�?W�����;��-�B�]�-�FB�0N����Ƌ�l�>�iP�^'�(U��)�JH2(VqP�^�����P�)�_'���(D`M�5��h�l��D.�l��B�O��n��S!<^֪�U��46����Ԧ^9�J��ԁɬU!g�d k*h&ވv�Q�7�D	����+
%��=�:v��%�y-k�0����6��ydDR�r�:�@tsd��g�4/\��Z�(�;�z��>�.�@�3Sl�����'FH)W�����j����g��d�J�_.]�o$� RƸ�-e_�[�䝹���>��^�^;3S	^�!C-�����lg���!er��m_�X;�mK���[a��y�&�P@��I�u�S��5�L��y�g���.����t`�o����0l}ǔuy���mc=i�q�Q����v75�'����M��$:��mD���|tu�1-�v��7�2#*��D��aZ>y���[��`��Y�}3Þ�y�	�V�UTv�?%cS@��\Nܛ�~�����(�I��³6�V䫐=�����h����|���I^9�zG����cv�vC-ƥ�J�� ���ֶ�����v�ެ�C\�+��WM;A�2��b<�vF��,���,r��梻�� ��H=+��mI�gċ6��#�g�2nJ���jz�����HH�y��")8'�Ϩ��4E�_�:)��k(25���4�y7�Š5`�3�w�X.����f#
��9�3�SqNgE��@.��� �#��cʹ�b�wvj�E��߼F.6�.2��^���C�`I�HFE(A�9^w�k���5G��'`K�V�Dl�4?�A,?$��G�~�'�=��b����m�TM����!)�F"%E/͢�/�؋��'ŀZa��q���?N��ܑ$��&UkS&u~d�I4��D�r=HD6�[��Xp1�[ ���������	iI�Qj�O�30_e�	(<��J*���G�fP��`%]��
<g�%�յK=����Ұ[�q��,�+�'{�_�%E��9C���:�GW6� n��R�m�;o���m��6o�+R��^AE{�N`qjx&-{QC���aoMtM=TiSxO[���+]O.���I�v8Î��� X��+M�[��ڲ�Q�%�����WO�����d��Ԓ�7ӒHV��,�C`8�y"��ο�Ԗ��՗�zp� �� ��í��[?�B� fg,"�cuN;���-?�R[���������ئ������`�l�#�PX*�Ӌ%�,6Ӊ���%B���9�C�Gg>�c��rg_�W����N�K��:LaR�T�ˀ�� ��U�>�4��D 8+c�(k#ۍ} ���4��M�����E[2+�)�A$�a�������IE�ֿ�� ��~���mX�ӪJ*B`*z������Zd��.3��C�{.�]"�&w�.B" �����w�־����墢|�c�*`XZ�Nw�Tg�x*��l�*f�R��� �TKbga�jX�B?(�G�X�����W�*F� d���f�b5M4��/h�~J�Ӻ��܃��N�\�[ϫ�ZW�tZ���XIǆ����T~�P�A��8u9���VN����rɳ~v���S9�I�k��xy��n;oO1�i�#���Pѿ|�s.�yJY�iI=8�i�c��:Rz�����t�0~�R!�3��/����'Zk:�T\��P�	�,���f�����_�TwX˳�k��(x�c^����G\�:X�IZ���N\ϫ�AO8��7	�8�}M�׹d��j:��!�cRG�>O�����vm~M�u�%�ȸVڤ�LV<O��Wo?6�� �}�6���t�Hp�!����֯K���˅GT����-'�X�/.ql��������l͸�ex��V�1��S������~�&+#kE:w��׀��lYx��*���(L�gn�����;ya�?�����M>5��>w��.�r ���g�stG0�J�L@6G6�y�Pn>Jc
����l+�e������GI�c�`%��wKվ��o�}��Ek1���������H��ӅB'CE��O̽C�\닭9kW��V%~^܊Sw����)3�\��H�W4*M�a�9�}�֪�f�_G�W�r4�(OăG�2�B�'��
2�����ai�B΂���:�V��ÿn"��w>#���㈇��u�8mm��u����"��>ڃ)���p��~�%��wD�ݨ���v� ���QS;�Y2�b�64-�0SW����{@7Zd�Op��)o�0���*tlWQ\��3k���e�bw��������#�@�gk���Z���a�
�6\m%I��J;�]�~����U3o�Mf��N�7�x)v�p�8XW|Q����}56�$"�'!�3sX
��k�Kf"��P.���,�>Ѩ|N��������u�zL���|�����U،x2��E�#&���%c�S�FC�gc�+L�t���k5�l��Z��f�����ˍ��<�j��k�Nr�ed���,;���<�e� P��n�e5\�-Nȣv?  m/����&��:�t�,����h�9��"�-�Hհ���銒J@Ol|2�=^�L@6ʅW7��ۡ��z���8P�ϒl%����r[�y ru{?���i8 �\��8Q��z+��s��E�����#GJ���5S��)/�O0�#o��k�̆�>����"�z���V�b'Ö���+����=4�@p
$Q�}���'�zU}S�uk�ợ|�J0��)e�Da�����<���r���~��q!5�]=�_0�%'�8���;X3R�5�2���$��d�׿4�B��:���K!>Vܼ�y�Hr�J�ɜ�Rк�i����.PJ�_�k�Ў�jՆCzDcWzq���a�E^�?,�����0D���X.��c/j-;�{��n�o���|>8?�B&��;	�݉z*��8jg�('X���}�x����|��w\IJ]��L��v����qoXk�v3\F#ZK
����������YpxG��Y���!��*��C딿��ŋ4:S0����<${�XE;���/��8���G:Q���LS%���h.0�y�V�f�Hd�%�!Wt��x�(a��4��a̭�|��q�!h�#[������Z�p'To|�^?��Eo�P��!��f�)�]����?c>6�u:8��ko۷{�"{9$b�y���c����j<�	��vE7�sk�z)�|N�7�1���<���� �k<_�7��^�c�+��o�6����7_�OOU�66D<�Cnq��溅;� ��|!\��ޝ�p��2	}b�����գ>�;b��ܬ��d�0�>�DE���t�9F����&{��u�g�(�+��}�>�Q��zP�'���uQ�[姂�˶����#�XPfw�4:�K���X粯���09�3���N��5���u���u(�7�b���%�8+G�(�N�2y�;�z��f�o%��F�|���RW�?+�j����MŰJlI�4s(�Gy�_j>��(��z�:^�wb�F���|��\�:-�c/��Kq�M���Z"�nU(�b�؜VѫY�&d����0�h��oņ�F��ƽ�z����+o
@� �"���0�����AnOkp�w$�nxb�i�|(]C/��<�jɸ�y���$X�A����4��!6o�^;e�}$�	��yRT~��A��>�5O��3Bw�'�jؓ���=/St�#�Ã�BLmx7��Q�P�ᠳ�X��pV�\\�N�N��oU��X���2p3����o1��~И�:d�����䁽&!?��S����dI�*^|痗�<�o�Fc����s����tp��2�n��q@�Y�<~b��^#j��Ƭdi\aiο�C�v�2yݼ}(Na�J
)2���rݍ>��Ӗ2a�Ǝ�q583���/�ƴ���f��Q�Ar�_��;Ҿ&8�x��"C�K�>=�����6��?3m?t�<o�t��_O	'0�M�i%��Ƹ��*�P���&-��7�i�)�K`�. �whv..o�i��P�*�z�ҖoI����[	�^��}C�|��46��q!�˿D�����o\�o�c:a4��K���P�.����8f_7��s}�u�_n�Bnh3��\��l�,J( �%lj�����y�e�{��&�<R$wG���0��[�ŇZ
��]|�0 ���,=E4E����:L���Q�'���R�K��8�$�[��t�����a,����Ac`H~��΢�����-Î������Ԋ�T�aW���.�r�b�ټ^й�]�q�Cxl�o���Y�W5^	��:G��.mf'�dӦ'Mwh1�	�����L���+}�ԏ��%Y�yf��-��W�y�0�m�Rf|[%����q��M���>Gg�o�Z�(��x�n6>�7�u����x�]����p.�2�C*{vf^�!�x{���`Kb+��&�5Ż�g���6s<W1=,U�'S�{P
 �qIR�qə�С_��h�yh�K������;���`�y:9"�R�g[s��Ӂ�q�قvo�s�%a����?�/��bQs�"G�'�Ӛ䷦����LL����{�'����2��,���k(՝W2�qKے_>L��Z3��cuV�	��I��b�~��џ��qw��_�$���[	�"��x�l��� M���������{M�<5�
�G"H����kɵ�[#���಍ 2$؆���G�)Z�U�Y���2�R�߬��G�52�y� �>a b
n�m��w��8i�7�'[���>��c+N��|��H�,�M���h��#:͌��%`��r52[������z}���ۈLáW��T,��LR�n�^91>�1��;�ʵ"K�d�E:�?��흀��0�kзB�G��OY�7.=0����b��ARX1��C�:�,�8�㻵z�����J�����4rG�+]��V��fE�+�/����'Z*������ܻ�wÌ���k݊���B�v63.�>��7q�ԡL��30�w6u��_Լa����a/oL�|L!mJ#���%���(}�~)�����G(�GjE� �˦m	b�P���6ݽ?+G���2,������x��&�l��Ry��>�/��V�~���\�*{�]�^W:Ӽ��a��)'g>��z:x��V��[Zt��wݐ��U8��ŷ�I�K�f��s��%=�NqC|�ү�L�_�q����k�����;��OQ��ĭ'U���O�m�7LN���uh�X54�T6O�����(B���bl���B��%	U�x�5��Fj�0k��O{��SD4�bq(Z��^ᏧPۚ.ox3Q��稜1O�;����j��Q�!�.g9��G�K�`�u"	NX��%�:mT��FC�0_+ (l�S�l� �q�8$
o/x�b��E�k��y�A9�p���{;�L��A{���Gn*�����¼��7�>u�u�^`�?~�mA?�/3;4��	4���t`n�
>��z���ܖ��X�D��r.�8>��,����Z1����װ���wA4Rց�N�y��0Spf���^m�~/��+]6��R��!��������&&�x���':�S����Jz⤩h!��H۝͗0F��j�-D�rQJ�L>�m �7&��*Ιo��4��ER7`;��d �:Z�)��E֤esjf���9����'6�gAy���a�1W��I��"�(�T`0E��s�n|�� �7��2�:��7@��o=?�3j�+R ���aKm� Cï�w�}lL���#?u;<�U��@��M++����U�e�#C�JhbɄ��+3�h��[,��/���T�Z��M�C��M�n��5�?)�}��>�%�%ܧ��'+����u�F�7�:�F�L�!�RkW�5J{ipç�!��)�~�c�`��S�&�He�ϯ��w�m0�c�jvk�?�<�@�h҈��À�B6�O9>� ����x"�`qx��@���9�!��1�p3���GjZu���L5��}�������%Y�sP���-Cح��H(bMYu��t��m��)d"x��c�"��ɸA*Q᧘��%��61�;��]�5�	����H�T�[Հ3:Kc�����8������\W�D,�=t|�|1?9%�9����_A�W^�&�G�E��⠦o�x�s�{,�����4��D����ϥ��>�R�M�O{ej���g�������ߛ�H����[1�!�B
!6E����
Ǆ��2�7����Xt3��a�r���$�b����m�z��R�d�~v|���P���q����&��1K�[77��]��@59����+���o�D�J�s)*?��>)��s1���\�m�S��=~�t�s��1~� ;3!��ȶ"O/֮� �0��fy{^>�?u2&�K��j���or5�fe���o���o¾�mQN�k�E��[g%����Y�*:�*zf\�]�F;m9��n���(�F4���'J�Eˊ�w�V1��B��$�Q}��E�OVR��	jV���z�%�������^�U
����8ow��K�
���erLu��Cͅ��`]1�,<ʉ���U��4��s��S��ib�P��c�?`���4�7��âw3BL6�?|���-U*�m.�����mR�ߝ~�[���c�b��-�8Ƥ)�4�*�mk:kX[��g7�#�@|m����ބ�	��b2NHs�|�'ޘ�� 'k4���(A�t��1��<�y���V�T|d✙.9j�kH0?�^�m��i@�������|�ÉЋ�@�ef�U�r3o�!UhZх$�		��{�>����єl�2U�1�B5%ck���a�6�
*Y������5�\(��fh�� 
=0ƨ%�,���6@�2$�XB}�~5�
��p��^�6���|i�� �<ć���?BU2�?��:�����&ڵ5�p,�C�.g��z�����R㈾&�M��)}�x���bt)� �(E�xEM�rE`�;Z2�8[�-*��v����H�d���v�}�܅�P�CW�'�4�����X����"x��.R����^uG�v@�5 *{�!� ��	��F�4���w��B?�k�p��9r���AB�=�ƴof]g�b0�oJ@�/j}������*H���}2ED�1���j��+����=��rK]�u�ˑS��1~i��۳�ɵ��M��%�|/�����4�?�邂x�.�r苳����3zjCk��� ��qߓG�T�o�	&��&�F�:��w�Zos��ܜ�+�Zi�~�Q��@��ƅ�7g���
�`P"��=~��Qt��c.���{֭.��;=�|c��`��-:4C_����)�G�DR9lE�v��sC>�U�Ncb�~|�����\��D�/�}�L�J��$�\��W�%n�_���`�X1̿�T��ΘT��	�i0-ޝJ���$�Էd�����sp�Y�0���W���md����y�m?�c W�a�%J�/x\W�AW�L��S�stq����S�1u��?R�����F8��bLP�w���O�x�/��|ñ1,y�zz�E��\�o�ߔ+��������ά��z'C�.����i�>#�}0���&�x�!En��H{��E���~z`�$��V9^6\b�	�#Se�N�C�B�g��hL@E�*�\�Z�w�w�ݗ.W�#y���l��Fc��G��&��I�;^���U���cύK����N��U�<ĜW}p[�:�t�X��l��5�q�Ӂ&�m\���|��� �-��t���JkOA�\�������)3����,�G֮l���2��������X��
��vgPj�^�|�U ��]�|�I3[����ZK��1�,�D}��n_��c>�T�y��tY��`�&������p{��+�햎6×�F1�|@�zχW�+�ȊW�����7�,�b/ƌ�����(g���#�ڧ�"��])���.Ҳl��{ �}�sy0
ԹѬ��[tqېq��W�p�zn\�J,�m�"$j!��}i�?����9�a�t�̡�7E����z�/��>.�A0����N��ț�8Vf�B���NX���WC�s��8�t�~������1��~�/@l��C�I�����(8�)7E�ju�w��+�6^MY�\ÈCS8rWD��'��̥��*{R9}��ٹ��y<˂��Rt��pO��"4���܂����-�����R����MI��뿨��f?�j���l1t����|s�w�	P#��T ��v�

��V6>�
^��BP=���i���v�&,�9 �ܲ�lC!���<��Xh7k}C� z�ܙ�[%�d�隂ɔ��0"��'Ÿ���>C�հ����[$���۟,���ö�]��� h0��#���^���e ْq%�=-��)��F�:�0���#���K�� =y���J��X[rTq�=<.B~�[٫�X��cf��0��̳�IJ\��	�}?�S����6!�Q뤌Ϡ���O����=�*0�mw̨�Ö����O�ͮ	$F 	��G�
	��Isf�����Zi,OL0&�|���G���`�rō'����2��I��HB	�{�o/W?�N����Bt������g�rך�c�W��'lL_�4��~k�wvU�������d
�ۤ��A��HnR�v�K���4'�ր�5J�a�3{�i���./�L(��>�n�{ͽo��o�N���ؙ����s�bv]Ao=�y��VD��r��1�#n1�j���3�܃�:$R��/�=�J\�:���(���X�W���0�[��tF�Ь+��ܺt�C:�ѡ_�*w���AL�
� v?��r˟߼�)za6:�F|BG20|����m&<��ۆ��m_`������x�X�1�յ��VT'�`�mʼ�om-�����PCA`Ǎ�L\H����J���7��Q�����K�n�l���S�"���Z���Ry�NUF2P���D�6(g��v���7Y׽;0��ӯ�(ϯXE��K���f�ʠZ�q�3�r����qN�t��Z���ڙk"��`s����Z���c�/LP�ק�%�w2`F#c7Tf�QΡ�y��p띫5x	
/
J�a�Xm��<#�G�C�A�6�l�֑ҧD7�Mst&���(@��5�.��q,Sp��9q�i/�Q�N S�cA�!7��Jl�/)��w�r�R.�@h\�޷�}�����oc�е5�*I\.�u�ŏ��x�^glt��qKN�#1e���	�G;����-'��`q�j��ض�-�_m��D��yQX�Jw���c͕��H���D��ry���@�3%b�`�P8$`�u)��z^�������S�\����y�������okO!��+ ~��3`6����t��>ۘ���z =gv��Vv���T��Y-ݡc����|���&����q�Ѷ�K��|�����I$�=�bi^�o��@���7[������P_TX��U�V�3M�Y;~�S�+����%O����V�h���ۿ��i�6U�A���c�h�jL�ŝ9%���d$�{���l	i�0��З�b�Zt��Y�5:��J�����O9g�;C��kE9���@��$��֧I�ճ�o�̈2U����_Mr���10�q�條W�z3V�]L��RΧ�_�]�� hP�E��U���Þ��︌�~A�����.K�#n���nq�r���e���e�}�s����g�h4@�QEޯFW��r�Mi��u��^����`͓��+�W�0����NJ��Ӂ����^�i�3���@�����x��/¶J:ؠ���Gׁ�"��
0����F�$b�3b���W����d@�b���b�@�_9۰��ӛ��>���5`J��et���KA�;��pcz�Ĉ�G�l&��[�oE�t��e��������o���Xs���d�� eW_s�v����{n՝����g�K����j���0��R�`͏{z(y7�����v���]<6���0W �BP���B�;����y:��ڵ�C牤��x�;�.��m�6P^M�A�sd-�m=�Ur!s`$O}��Վ?R;����P��5oLNNʴ6�{�N%�G~�bz�K�������c^�5ܟ^zo���yR���[��\J���7����� Q (������cjDl�A���"f.G'��(�%�Q��z<�X�:�Ry�|�8��F�V��h��F��&a��;�f�5�)	�{ő�"Yl-�J�c�{���?3,� �:�ڭ�i��*r�[>�e�B�e�7
�Iԗ�'Z�O\rO�p��T�m�5���v�Ci']iR�Idx�Bnƺ�c|��	�Rø ����}�/��n��� #���|���g�iL�� �՘��GL��`���ob��4��0,��>�_gnɌ������*/E�y�l�3�#\\�UPȎ��t#�}�:��\v��D>��KM}�s���h_q���7�7�j�v\9�I~*���\�I�{t�H!�t|�ޓ� IHԌI��{�z��5
�P��\�TMi&�h ��=�D�}���)ȑ� � P��V��0 ��%����볭^.�(���U	�#��6g�sd)�#��D�[� �#=:�k��eL��ˡL���ߏ��+�"]�`Q!+��60\ptrb��o��,�шt2��ͥ}��@��[����pO+þ�e����lD�	�)����S^'��������Z6E#�Ǧ��j0�!�I�SQF�y�c<B���s��%�l��~�_�a�4j0�n�92#��������M̺A��Cy�k�����-U�iv䳃����� �#�Z&�z����!�~^���K�K�������>�ȧ��2f�8��b���wu�ɯ�����B>�	[^[�5�q��{��3d��@A=����?�٣hXA�^�:�vz�9t�o���s��+����ye} y&��\M�RI��du�ĭ�͜��Qs�j�H��;�Ml;Pa4y�������=89){����]xl��)"8�Qj�v���p�u �#���ܔ�p�jÊO�Q%�}p�N}s�_|p��QF������������a|.7���x��&m��4F�Pj�\*4�GDj{��X�#{o�SE�>�뫹�b�+پ<���s��_[��j�O�tR������=4w�,P�Z��)k���ŀ��d�) Ȝ%T]l��a�X�Kh(�ZL�>f%E�zª�&�7P@��9�o�IqJ���ۙ�<W���������ʃֱ�5��*-�JK?�8N�"?OĴN#u�	m�	����{C�^�z+�]P�A�9(CU�rjI=�E������;����Y���x��i��n�2)QXd-�:�����(`�q�t�Pڒ�"t+LѶ}�P�v�|����/�.�e���| pMK "�B�ډ�дuhm�v�Y�wI��������4�� ό5N�iBT�E�
��J"��c�3(�1N<z��gs�rவ"� wq��P��m��DH�N�d������u�%H��$��ϖ��S�pl�9��ly�yAl�?2��+	W_L�>Ѷ;Mulͫ��Q��U>����1C�����s��ل1����\bc�7�J��`�{���kڦ��e0f���i5h�ߐ�J]@ ��{c4�Ҡy�}ZZ�4@rA:�δW߈�v�2�^�E$A�Y��)�#�٭(����d���G11�Z[(�Uڨi�=�v{�B�҄�S�I�gv�N�vv��������QH�XOj��s� ��Y���˅ϟ�,*4�,!�� ����/��
X��k$����3z�E� ������-��7��j1|514�[� �m>GK�o�|~�Â, �hb�qC��TiF�i���a������R�� A̰ATk@�xE���_���ƄY�:�8pp���w�����y<ˍ�%��ͯ�a��o�-��K_7%��x��I�a߱:�
�8����Cr�5��0�S{Dǈ����?��d�8m�����]�i�
���V�ʹ})4�S����f\���JO���(!z0��t�;g���
��o�k���e����h���D�`x�e��η���wѺ
�S흆GIw�\��� g<�v���D5"��Jd�oU�jőB�\��"�U�<�kP�]<�C����C���'+w�g#�!�f6޶����� ��2V�8J��$ћ�-��T�cBŲBh�WĚqxu4��D�������)�:/9�����,P���p�L�W�ٰ�w7��Ez?	�;q����H��������:�����L��[I��N��*e	ܣ��?�2l���j� �4��5��;�ؐ4xM�f��u �3fO�L'�c��N�
��(Z�mm�i@��J�U����*�US݄/�J��bc�O&��P݅�T���Q�������:������i@}�dh�Op�b���w�j��.��>;��+.[�������6x�QtK���K��F��Y0ZaT�|�� �k�h�@�+�P���	vu��v8�keA�"lXT����.�(�̜��o���k��ӥ���n�˿��Vsϭ�W����Ii��J�7/;��5DN5�=^�7kz�6jn¹(��3��tHM?��P�o�=T�7���9+r�}�N�|�~3�����:)&�N|e�U�uQ��"���׮LD��.}����.�H7�U�5�k�E�����o}"~�̦e�Pm�S^���A�2`�d����=��{
}ٗ���:,��tc"Z��ع����������-�����(N�%� H���y�Eǁ|x@Њ�e? �%���eZG�Զ�(:d)#�!�ᶂO��"�w�!���B��!�pG�L�N)�Ou���M8��M	L��7�F��O��;��wǤGF�_����?�HN)�"+�6g������r��@���+,�\Ј���{i��0�X̐;#���;�g�X�L!�@��
��6?c���~	L���8����>�0�1��4|�,�Ha�c�\����ld�S;k?ʍq6s����,�Ҟj���嵒@g���aqI��`��X׀s��l�N���|��CPԀm��G&��Gye��/a�LE`����7S���0��L�g��GЖ\-p��٥�Ɲ��P|��f4\!.i�ҕe0~���A��cu�h�~��S_�X�/�XJ�E��U��L�߷q3�:F��*���y�x/2v�*�t�g��oDz�a�W��r�Z0+,����31�ިh��>h5sx��'siy.�sr���.\�KrwU_����� �t��:A�'c��Z�*o	ԥ�h`��
e\��aӴp D�|{�g@*~'��h�m��e�L�KR���a`EK�t_,`TR���0�|����N� �c�41�D<|Dw�LSk�ҭ�D8�bǂZ���q��j5GP��l<�@�~ڷz�������k�-��-�O����Mz/�or�����_bz�@Uro1u�;z�W����h�lu��3Ŷ���h��R�'�C`��D؇�}����5X>(񫇽:2�3�P���-�Q�S�
/�&��íJ�8ϱ�Q	����7nڂ���r$%��YLٮW��ő"�M�Ɉkqz��j�Y�=j�5�M���C��7!{v�`��Ġ��n#+GW�	t�m�}�2����N�}�#�)5[�5b������ E���!1�������œN�k�V��T�<L�o5CN��I���38%���UB�]Q�K��Τg�sD��o�t���-O�h�������W�^��V+<h�FW@��'���wT�lߓ�����m��d�{�n=�Ȋ����F���E�l����ڗS}���$��'��J��A*AŖ�W��I���l��@j�q�&���4�@���+KP���w�A^��5=��t�[�Xv�<�˟�,2�a8���q���p�{��47���z z��Xp%h ����;��5KE�AW���*ة�?����I�&@&�%��~���ى�4��.�?2�<z�-(R\�x�6���$}f��u�(*Y+O�Gxtzd{�,��=�\m� ��#V}+ʳ� ʹ�5��k5�d�sp�Ik}�c�NE�D�y�'|n��غ�����*R8#�{E��<�ؽ1�"Q�ݚ����[=�w�u'����\,q%�ӣUe�C'��r����̦���Q�r�z7W1!(��tcՃ,��F��e��Vz�G-J:��M4��;�Ue N��VN�B`��a �)~H&[�a�ͺ��ۤ�u������5�$y��kN��UqiL�:e�r�{�#��D,�/�֮]+�?r.�_4E?mU�&j{b������p�I�X���Fr�l_m�����o�Q�D�c�h�|���^�F6��U�Y=��۽�ѯ@ne5���� J@N�!D���e>۞�K�e&ݕO62��%T� :c��B:V�å��8{^��]�~!�L�Kx���2��ϧ��S�L�"�}�?T�$ '��:U�󐟺T��va�s��oͅ��R}���п�{b�A4d*q3,z�QDc�ZO�&��q�U�YMEm	��GD�v�5v�� ~[4)m��r��ѝ�ڍ6�q�g�4��}EEr�w�7������j�r[`y����e���	����M$���^���R�4T�`��u�[����L<cp�m.	j��R�@�1Pek&�����o�g�]b+�����䄯VC�#_���_���N�vo������v6�}�-�S�Q���?��)oq�&%�����M��̋W���r�֪#|���>R�m{~�f�ȖA��V��b��ü�U�Mi5b�鿈l(+Z�@q(y�'�#��Z�&0ǟ4���>��X�>�Vv�Z���K(�B�V�%D(q	���uW���l��p�˶�h�����q�E���ȼQW|R\N�x�r������Q��SZ�zC͂0{�M�mJډ�7��Ug_\ HGO����'߮�W]M����-��nC`�=!�?��W�Ey���9�\R��jc�7� �6\㾕���+�Y8j�6b8,6�ۜ���``0wt�~T�l�E,³dGn��?�94>l�Gu��3�yly8��mÃ��{���� a�%p�� �����P�������Jd��oR����s E�az�]:�z+�7�K��~�FF+�~�]C�A�C�(��\t�Q�n]�O+��'�b�q3d��M���������W��v��@7S���Y��/�._���H2��p	&1�hS�-�kHt��PmBՔ�8�ޭ�U��N��H� �$zu�Q�&2U#�b�Ǖ��E�K��])��9Ӝ'�=��z��$:���Jk�:�;\��TU`���f��U����v b��<�k,R.7�L�k��+1w��9�>D�9,�0#^i��7߅�����⢔cs�?H�D��\����| �p�G���a/��8�K�X�����<K���8�W�mT�GM��R]!}q��.��	j�����O��gL�5�3�b'E�-U��ǣ}B��#�`b
�u _�*��+3�-���m�ƒ�VM�)Z;݇��u}�T���Y���Vp��#/����)�?`���f��U	��F�.��%�酈���+pF��2t�*U.K{ɨr��P�k"c�"]��k3���l�וFi��-k�1�t��$��d��=m��-���ϱǜ�Kb����X���|:^ֹ��V.C�&��N,������/�hAȎ�<�M���u�����ߙ�8b���{=�H�:8��K�)�쓢T��j*s��O#��&�M�cK�ȗ�������9�3_�G�E��/�Ӧ�E��"=�$Ae"Y�^(�ޝ�D%0_ڊb�9s��1�"�S�q�>Yt�)aO˭�Wp�����r=���9:U����Q��:��z�MJ�^�j�DPa��H��YEPћ�zW_t9�q-���yt.�i��L�43��%g��6ž�s�;�������S�1}��t<$P��?��~|�&k3R�#�r!K��B6�Y`9k΀�i��Q�� ��³-Y�˅-��!�i����,qd~��;��f����9gÀ��k�?5�#�NS0�^�#	��_�Iy�q4EAJ�4�<�#/T$�!�y]��� i(ĺFһ����T�����C�H�.v�Za?MU�ƪ�KZ���H���b��v�:�L�٬q�4������XK%by�w�d�Tk�Ȥ~�r[j�,G	���3k��_n��=�#u�9|&�d�\*��[#��n$uϒxHk�ȵ�^R��4�._�Y�aFUU�t��'�����f�Ȃ��_Ў� �>��!��@�����z��b�U�ܛ�U���S[�/��NU��4��5�rnu� �!�r�-Q�	��̇�$C�M}'~s��n^�����WJ��ie)H�W%E/��Bu�+ ���d?Lc��&���g����>�b����	�z�@�u����n�(g���0�,C�"���U	U=�9�}%����x�@�Kü����TX�%u�9^:FW���E����G��W.����,�uԤ¢OJNNwD�_��N���)�\��h_��@Mo�`���@��FM���[��
<��1�<L�zl'D����:�_'�|\&��V��VB ��'I����"Gۮ9-:<�ej�D$���T9	�.k���䘂i��Յ���w��^��q������ޖ,���M�U���Q�����|���,���)�?���\�qB�e%�6�{��Z����ow�`�U����ӍF@U7h}bv��p�l3P�I(3ɽ�\�����h��g  H�����B_��xFU[W�~L�hDOk։�Z'��y���v_۱;�2��� r��N� ��2Ȍ�$]o��Շ̉��6��q/ć�o�$�Q��I�;�i��(��;j��%��f���Q�u� c��M��=���4h�lq�{������ C~�U%�8���/��ͽX�Tw]ނ��G�hs9�C,��x-�̗Vjxq� 0q�
��ri2=�u3O���^�DP����M�s$U����>���n��0��S��c߯�����JY��T��Y*+���B�\�}��y��>O�����-mx�n1E4���F��H9��>���C���Z�ݢ��Z8�h�.��W��W'����ޥ?+n��+���G�h�i��� �9D�B �< �szGQ	�������H0��9��`�w*�<�h\0�^��nj#"�~�������;�X9�A���5��1�J�|һ.���[:�Z[CTz�k���US� ��L}�Tҭ�n|��fAG�V
��>{��� i�P쀁O��]I�u?ӌ�R�49u�{yo��ۜH$�*��	p�M	2G�SX��v�l����C#e�j��+q%�gX����:!M�5Lr�j�Ȱ���OB���'oL ��<�� �M݄�h�
\�׋�*a��~0pX��x�SP�Ph�k
�*En��XPe�_{��9y�A|��$�>!�/�2�����Qv�7���]ԡ`�d�,�E��e
���\+rZ8�˃�`Icn��iQE5F'		>+�I����ٿoR��ȒG�$��`��6��������^<B2� +��b�6u҅r[a�L�y�Is�&K��fβD�R�,�؜M��k���,Ǝ�h��}�Ż%����ɽP�]V�:kh���i]1��?�i��<����l��{� ��^	/������2b�΄�a�wL���2���>�_��Իx�y'� ������g+Ѯ��I��t�;xR�U ����"e��b�M�>eF�5���,�&cP/&����9+�Q�@�6J[�x����dWln`�v8/S����f��n\�!����=e����̘�?P{b��{�V����`�=d㜖έ�"��j�q��H�Ԯ�X��\�pqRޛֽ� $,O��0G�ob'�>��|Q�s�MR3�h`�mK��[���h>�}�Liѿ!����A)���!�C�낦Q� 7F�)Mas�A*�I�x��t���8����A�D�/���Ӻ�q��3�g<)�Ŝ�g�Q���O�Wk��m
N�G;dͻ\���[��3�����P+ղ�l_8���T��9��J!u4��@�Y`ɋ'��_vD���̍H�q0�Vn�Y��2�m�s$�#��:�,8���U���[�}�� �󷰱�����h�,���2�U7�xk���B��n�O�4�B��ov�O�g0Y"��A��@�RQ̿C��]�!��HL)ֻt�mC(I�T��x�цk�|�}6��(��9U��.���D�2h���j�C~A-���JЋ��5�T�u�.%�7s��P�ǃ����9z�Q�ܨ8�rg�=L��O���!-궇#�n?�M�#�m3����������짛A�p.pF�kK�Y!�H�&�MY_���e�-i`!ϟ�UM{۹Z�Q:�Q�rt-n�i(�9�j�����~��b)�HHT	Ü=�lSv��������z�2�[���q��A�����^t�X�,ȍA��*`�Ĵ#o�=$�XJ\��ŏ��dz���)} ���4��FT�(͓H��X'7s����(��"�4([�p��D��{~�Y�xr���Fx�J��'	#��ƪJ���<�O7��@�7m�c�~	xl3���19.��5Y)� ]��%�v�JEC�*��:	NF�U"���ZVQ�#rS<}DVC^��Jjr���a��H�3֢���l�y�3��B��,1��0����n��0M!�p�q�Aw��\�!��%�Ê�����#(��E��մ+r�����[Zd���xWkх����&���Kי'�pq��G�Hϩ����<I��f�]�{8[�PU':<�cj��?��="�!ڹ5�u������N`�:ڳ�HM�X>����S#&�rV(b����X�z�OA�ҫj!4��^��
�Rf>n�'ۑ���%,+^%���{UA]�g� ��0W5���Rk}t���G��;!�(=���_���K�B�֨#��p����޶漠9���N4J�į{�J+�6s�g�=���!�S��~ z;�܋���C)#�ZS���[���[��Q�ɶ�'dK(�a�~�,D����~�"��ب�v̔�O\p|q�S u�5�������&��LϘ�Xw�`��xM^��*K5k�Q�c,c��_S��9;$-S�`JA��l�C��C7��Ə����>�|-�a�P���%�ʌ�xs2޸ȶ}�x�Z�,q��5D��	��)ŘDQ0tMD�����Ỳǭ��ȣ��4V���-|5]�-�,U`��&���E�O�; �z��5c����A�qҭ�>�0.�\�$^���M�,�m�M��@
1�#xU2!c.h�㭓+���;<�nɧ�漗Җ�������q݇מ�\W�;m�#қ�M�#BkNo�
E��<:̨�:���7;��w�}��~��0�Q�1"�;�9������4��C��DyZ۾��ܪa�Q6��0�������΢�W�UY\}퇃��M�m�.~n`W�\6r���zԼ�ӝ�\�W�в���=�b�s��5ik�)b�Z5Rxƺ��#֨�|�
�r,��N ��u.��[C P[
a<�4'��4(���3�T�^A0oC_4�ɭ�V������=ނ�9���L���Ҽ��WKE�8O<��08Z�ni����5tK�gj�?ghd�LC�~\,�́��%�5��ʗ��6tz�� ��h/�]x���+�gk^�%I��4 I��]'�����E���ʽl郞���Y�:�]�X��7%����1�@�iR_���ؕ\_C�V���oq�~�D��e ?6��,��Κ�Fl��*��;����I�Xp<s�ߜH��Y"�ٸzJw]�p��:���-����a��N�c�2�Y���fH�'�j�:��o��e�֝�yDp�*mͣ񅸅�,v��St>���Pѯ�]`��=��RuJC&�����?�zt��L9��%��;��m���%}��d�`@�_���(�T_�� B3j��њ�|�^e�\�v"G�F.�0����$n���oWx���`��>xP�:emڈ٘~��k������gJ
�����Oz;q�Ƌ�9%u\��s�<X*G1���m�A�	��C���&ӻ\�L��d�>�F9^�ȵQ̞�ʭiIm��n�V�\OJ+�"N�
t���
h��p}F�i�g�S�c�l:����n��@3!�K�v� �p{���ʆh�����vP*y�
�#$B�j�Ј)�"o�7{�y��yT�{3�5�Oa��\c��X���*�/H�[M��a�eNÉ��V��Aȇ1SF�3X�$�/�٧|N䙫T�����~[���ْ᭰�6 X)~s��N�Q��ԩ�kzSK���3��9[bA��O��y�3��	����;���^��Tq�0$II��v��d���+�9�4�؛  ���$��:�G#���G`��π>�Z�Mo��Y��Bk(	�gq�˳�nf��cnA���H@�Mϡ�J�tЯ�и}���f��[\��X�2c�UM���Ťi���0T��3X=bQ���g	H�� ,�N?B9�s{&���*�#�m���#�D\(G��T�R��w���vg�'d�R�=�~|z*������c���)��M�B�`��o����\;�=c渣��7y��o���g�=�;��l��D�Ab��{�d��C):Z���P��Z�N$K_�3�ET�7U�����
��D�O�feP����)�H�!kK(�ľ��I>�o�8ZH�%����yK3���۱\LZn��V��5�]P{ o����P�Y�ț�5�Fů[��3'�|�.ZB.���")�SiLޓ�=�p,�XD}n!)���?;�UTW[W<�K�vR_��LZ�s�܂�%���cA�D��k�3߮��f�[�,��n���Щ��Z���1%pe��_�����)��Xw�'��t�L�������17���Th���n��� �ţ���9�H��)�'@�E"��٥0�+���r��4r�3X��Q�+�FH�u��!�7��/^)���+{ћ�EK��F�k�?k�U3q!앉_��5��c��br({RY�y<y�oqI  ,���v'>�)��6|cxw
��)�AGڜI��\'������ ��jǘ��5��fa�����V����|$s��6J�}���o��'���^� �����0LqbfrK��az;<���:x��sa�O}M���-��G�"�vv>(��frU�_n�#�!��Ph�4��?7��sk���k�Xz�f��6J�,�O)�>)�Y��QZ�ҫ(Sxw�/�7Z{��g(7դn/�<2Gz EqI�o�h��R��6uzP��	-��z��y�M�����iU��	Cf=�cdN�Σ䍧�Х��#��]٢u�#�J2�rTG�U�Ӗ��s�9��%�_�[0OZ��B	�N�Fq�昪����k���>x�cWL54�HG�\&X���~U֌�n���m��%��z�{`s��}{JT�
�;�j�累읿�X9�:#��1�?�:�"����C`�"���H�7���}�����ś��U�ʎ`���j���fL)F���:WX8Y�^��"����n�=zL�Qh�� _^x�xݽ�`�l�����<���V,�D.��������,��ԛ���C�a�n�R��;� P}ǁ��&G�-�"�f]�Y����K�ޢ��->sbt�RM%.��O��tӻ!�l����pDiV�Dл`R$���o�Hn���8�Z?C���!>Lz����$�̸�xAБ<^�*�:�)CV��r���*�Y���������r��*�6E�P�F�|���E.�z��y��D�ϑV���V��+���x/���^Fh�Ldж4x�N��my��9����{�w���i�d2�ҭ�UPZό5U�Ak֙��U������~���I��<�}���lYS¸�/�)}d%ڪЀ�W�zޞUAd���S=�̟f�%H��89;!h����? 0b�,�.�Y��MF0��������x$���!�>���s&�����&B���)slA���3G����E��D�3��]1xׅv�b�c+��AX�W4!<3��~���^ET���s8��x���U�Tg�A��~$ ͵�=E����D�U�l���ڢ�N�H�D��M�<��kmj
ɱ�֦����lvP�ˏ�7����n��#���C����V�a��Н�HC�U�
�{��(����c���Ty�_v���R/k�amOS ��w.�8����oLq�CW���m�!�$�� ��5Ǹ�Q`ѳu?�������W��-��R���f�?��J��/�<<��7�%s�U(M/`�ɕ����O��,I�OŐL�:�q.&���lq9[-�O��	��}�3H���ͬ�]��F*��ts�'���B�$�j�c�zr�j�)MU�~{���BRt������)���9��,��e�~��{̯`ۢǞ���*o��l ���M�2�����H���+�8k�
�# C�:��յZ>qUZ�� ��_G��: ����YP�m4B��ﾗ-�1V�����F4�L ��v�̼}q�������xN-���<�m�Y��>z7�J�E�M����xQ�!e�VV��Z�$;��3�r���@uX�[��:zKk{�6�Y"����L�$X�쐲�-5�{$��~�� ��JLX�.�Z�J�Z����ߐ����������~o; �&8D}g5�������V �;��(WeO�q�:Qe��le�c�uP�o�Έ��uS#��3�/܆���c Љ7Ӕ���N�����!�ʄ::�ɛU��\�-�����ɹ�����J�$[���8)�l�'�i<%s9_�^,�h�e)���Rr�'����僚ȶ��Z����e�rcvzY�����!|������~Nࣚ��+�*0��?+6�%�d���`�w��F������LZ[����-B����@���n���Y$2`4���"���N@mO�=̖���M,�r�1s;�,PΖAL�8�%,����:	�4o2�y�tuN�$'�wj$,������a�9�>�N�k��=����̞U���c��R���*�	ue��=xSʑ�T��`��Ɖ�G��O�Yo�"�sy���`�)�L��18�e��Jʮ��_T�{�1����=\���&n2�֞�mn��F��R����/���U
�(���!� '��d��XmW7�_�B�y��g�~�aR���8��Z�f#?�w�1������Y����΢�|��s��Y-�a`R���!����@,B�>������03��(Ñ#�3�v�B�l��g�N���.ɠP'�GEM�J���Ft<VE�Xs/L�D�4�����-��[��:��CTZP�r������[���|'�y<�T�	���F}���A��w8�P�PFFeb1
�X�|��Z�_��bV:�?"ܑ���8�9U��@��"�"�zp����J|�1e �_�*�lǢ�>+�NP�[��4��Kli���ύ�3�lz�S"N$ޗ
(�1��y����><а�����p���r���ӎs�jC��Cx��<O�h�*�E��#:���s5O#��Hh?qGy�hx6u�A���bX�x�j���������,�].��}�rX_p)���c*�J�V�c�VsMP�b���&�"(�^�B.k��f��U]#u���n�Ӎ���v�܌|��hws��E}un�X4\����F҈_}y�G@=���3f^�y#��߈~;\���@�v�� ~QN��?���C�?��
vo���r�M"a@���#L���� �")t|s�}�՘3�T�3��@�Ԥ�����O�%�>~��Z�)a���^��M�e��@+p
��vZ�~9��T�Jl�ypC����
����[u�x8rt;�p%rIGd�C��SjwA��DET"X��{�[��j�3������;��"���ʮ������̕+�Y�UH7p�"�P�|�iD��&7�������"�����x;��瀣�jH��(�/T�<Z.�M�k��_����sv���tr�U��W[�Gl�At���gP뼿8����������~.��ՐG��j�SU\R�P���o������:�O��Aj�ȂA1ɩo�������-�ie3����̬3��U.W��bM�H�k9��A�WD�o�s��Y-Z�}���ɫ�w������� >;g�9�c)Jk*�:��.J���\�}GK��V��� 9��bR/>p�����'���}�XL߁����9�h^u$����߰O��Rt;H*�g$�/(��N���A��̭Pa&�YǎF��@,���pV���:�x�˃�Z�`����p�ɜa�#���r��=��ܖ�U��W�PHɟ5��-��+��;��_��k������)}��L�Z�Γ��T2�G�̈́_�/4����Z��!I���;�kf�~��y���CU�zmwϤi!t��w)*���K]��p�MH�==��VQ{�i>�>&U���`��K�O��ᣝVE)�֜G,���xu�I��ɝ)j��f'2=d^h���B���~������{�R�}PQ��&���,K����� ����^_�:I>$�X4�,���kc�g;���x��/Ȯ+7F�g
NE��8�z&*�]�h����T�t��p��ǿ�k����E�ǿ!�g�z�������r+�H��8ذ���{�X����B�#n
j��/ԛ�~�=��d�0b�����Rib֟�����������H���sweDZgE���	.��f����x�\�b��Z��
��o�S���g�����V�p:��g��r[>xo�7;(U�Nr���#M��	�B�~�.��?������&�׿8��UդW�N�M%�OA������@��(+�9w1k����Z�;���i���p�`z^E�>P�,;kx�kNH��I��k�#ýFe��ʚ4^��^9<����e{JɍP���7�*����받lc�]�W-���lƍ�G,�D�|@i5�&�y0��;�"�T�1���R���$|ʘ�I�/��pxϽ�� M�OlS4��s�G�G�">�|�_b�'��S<Yr�S\rˍl0��R�v��a-h�����J�L)��əעS \0���~�s��<^a�H�<h5j���zcG�H�5�X�}��}Mk�W^��#�!B� �'A��q�� %��O��m�s�1��~��Z��US���K=�vvU��w�[(���8�D��Bm� j�X�Yg�p+_!�D�$WSu�Ǹbe���[@��m��/\?�����>�k�vH����g��׀�{7�a�ƚUK�i����DBi) �Pq��@\[��JL��������E?��v~OB��I�uZ?.H@Z���o�2�mJ4�&����1���ۈF�y���6��z�}Z�]�c��tL0fm˨�>@��O:���֓�#�3��V�xgZ�+�EW�s!��4-Q�,��ω.�rm�#->^���0�u&��XRJ͛��L�4-��pV�7�bG�؎
��Q�D鐵w?��BXq�P�;��D.:�jx���"��]F�v������0�k��6L��ml���� � �m���/�[��n���;���c܁�ʵǘ�4BK.x��%�������@d��K�X[���f"O�.g�Ev�D��<j8�o�CU
jaL�nvp�ޔP2�˖9TH']5��\�D������2��oӅ*�#o�G�a?��\�����R<�]0giN@␘dӲ��z��0�Q����T�4�8���S36��Z���A�>ǵH�T� ���;A��-0�ّd2У���6(:��T�3�i�z�)k�`c�W'VUl�M�[龃��U��su�½��M�b$������-/��3�޲?7��D���m���Ҍ�\��؃t���n6�$�d��ӓ6����_ܶu�܊�M��6��3��g�U��f�Q���%�8~_\�а�����T�u/jS��:��^��`���nY���֖�ALg�W���Z86�̢#�Z"�M����;� ��M�(T��G��`XPүBǄO't�2��t{*"�������z�z��I�Ѹ��ƅr�9L`��H�h-�[�~�frK�Fgs��U"�JC޳��V��]tYo��޻�zV?�j����;��Z;g	އ4��P�I��Y߾S��H��6!0�1��{�;��E�Np����TtZޞ~�=L�f��0�TP�Cٴ��Yke�� ?$&i��a�?fxTg���E)��R*�<��J���x���$�z�Y�+FU^�,�Ǉ��dk��~�mN��iuآP�,h����͐�Kd�3��]Κ�t��8�S��QtKMdw䅝��4�k�t2=�yE�9�S������w�8R*[Z"㦗�W���REڠ�h�<�=O��H�k���g�J	d�-r�P�s Ыd�z�M�{��I����ڡ������Ԉ"��	�r�k�݌�%�&����y��,�ղ����+z�Ǽ<�>�O��������ߜ�k:�4	�}�@���b�Ҥ9K�9�X,�*�}���Do�_�T��.+�L>�|v�5�K�Cv��BV��)q����*�pet�FU�Tn�ɉ6���{�.�h���$�i�,x�@^K�}���}���5�D(�o����Bn�$&_4g$mI:�Z�H�FY��Due�Ư����sʛ��q�e��d�ed���YO��28J�N�2����ڠD�k�XG,+䂥�^zh�����g#�P�L���;��:B�GrBX���)竷��2��)��>k�@I!�Z8~h�p���cf_6��ۥ��T�L�6Pv���=�-��f{F�(��M<��3j�<�K��T��+8}�����<���/�t�Uא�g��Gj>G9,�{r�i�	����>��&�I�e1�?C�wג`,��V�2�4����t��#[!ۍ����V��*�����Ӱ7\x�������N�.1%U�Q:=s	v�֜1��CUS�a�g9���c����s��z��)����S�kGH�Y1��n�m ���d�~��=������(i���Ƭ���PӀ� f]��ʼ/Xo��;p�k]�1PG�������?`D�%1^���nD��T�N�.
��z�䗗���Ů/5A�ϳܺ��%=?r��Y����ө���,Ǭ�%�5���1�U+IyZZА'��
������#	_�	���c�CQ�{a���B��n�MøX�ԧ���E;�C²h���
7'��Ve�^6x����1W�ɕ��ȴ'���4͔.<�~Cs*�͏�ԂHܷ:]�4ڹV�y��m�<��:V:�j)$��p(����9�w1.l*n��M��I\ ��ĸJq�沗2b�P�6��`�7?%��<"eV��4���P� �IY^�I%Y���AS�0�Q�5k�Hh�r��["�5ϢM��P3gvxTX?m���G�ym�+ا*vE�C�Ι���1Us"��`U3u�ӛ6�L�_,`%a�rI�*6֝'��U�TR<����{�E��%��p�K����������-RE���.τF�ݫ����+4v`���~�X����}G aN^aqH �$C{!�3�%���l[t�;i��%k����3^�5��˽J7{�u��X$�R�)���h��<�{Y7�w&�2�@�r�^���%a�\�mWsr�۬�eV��kLr�G05�ܭ�~9
�LJ���0c�ix�߿����R�J�9�y=����)��|���<~�`��D8"�,_�Y�0�QŐ����(����\�� �*ds�&�7��$������*�tǓ�8��|�P{�&��C��Frf�+��{�����g0�^��>��I�rF1e�d���3; ���	hޑ��=�+�d)�N�*��H��)��zZ��bB�w}E���u0,�������Cvu�2��Ȧ��>���kZI�b��9��1�y�NQ����&L	�$l+��w�<ԉ�t�DP�c!îG���/ WbБ��!�S��V�^����|T�b�|�=� ڤ��v��b��1l*�A� ���u�]���F��˜_���t�c�Dq�-]��_]Do� �Ѯ�υ�p�9�fW. �pbp�p.��.<՗].�	���YXr�*v����,�A1�L9^�0����z`��*���@�f��x@><Y:�J�R�F�:_��y>�w�"�`���"�6���&�������i�c�b��[/$ C�ek0M�t��Y?��]Z��T'��C����IK�
"7��5��?�e$�+g!�"��"_U:��N.:�;�cAəM��N�9�f֟�P�~1���*��恄n�dm����;�x�5i�-L�]A�]��� �t��k�s$|��[H�����}�1�Ѿ|~��?,e��JB�^Ң����z4�r�vD��gɀ��f�y'���K��qW�h�4�Y�HR�S�-`Pb��X��XE���2�L42m;Q�ˎ��dW��CW��1��ta�ݛ�����`��羨�� QZ�c�Q3�P%Z�%�������|��q�{ˇn�
��0����՞�3�2�b��{<|ԑW3�ߗO���g��'܈��ɗ���~�SѷG8��SX<m6�:�>�I��A�Q�|~V����i�W��~��Ay&|a��
����*��-��
j�z�!��m@iΜu}+�p�H��Vo�Z�R|��4�|�AX`���P�b���Ȗ�~5�^7i>x� ���f+����7P9sw>3ψ�c� m��c@�u�<��F�Y5l������Q݃��ꕆ]L�F��,��bn�'��)}���0V�Z�ݞ���aj�CE)��S��R�S#z��Y-�K}��6��W�vۜyy��D�n��QE��+'��8�U-䱠f>��St ��Y��	�c������$Rj��^2�Ʊ<�=���B��ٸw�zˆ<W�?bnRl�)���O���V�;f�Z9���7|
+�@�+i�2�R���A����I���΃
�&+u.f�hI^p�k��疼y�����F��2�#��?!��^�}���G��T��B]��h]�u�����0�is�+�����w��.�1��U��s��x���U_��b��D��$�G��l���Gc;��u�c����z޽��tה��1�ΗQ|L�S��_	=D|�tɷ��h#E���?�&S�����s"HD���5Ճ���ns{y$<�eZ���e����nRh�����K�>ܔ�3\�yGo6Nq�7T|:B�Ύ�N$_J�j��aB�t���?<��f�n ϋ�)vG3u�auI�=��C����4�{76��KE?}��ى�c�ې��%
녉�Bƽ�u�����r>�E�}4
�T�)F[m�=�T�x���V��������Q���pqaJ�S��<��y"5`$��9*m�;<��x�k�D �PϢc���rQ��W,tK �����^X���i�ʇD�f�kq���:��n`�)@.��~�Wl~X�2[��k��S��$̄#;=�"�#&����R���n����m:R��qP��-E��Ė�������1���&0��L��Tf�~aŀ N�������Ȳ�o��c�
�-cl<�yf�p÷2F���]��C�Xr`I�!jX�3Y[\v�Q"�O�	5����U�kU-��gA1�%^�ה��<���o�?f�[i>��?:�I�x`5Ƨ'� -���&�润 ���9��)�c'Y��v�� �S��kSm!���
L��^@2z�f����YÜ�]�b�>�^�(���f~Ʀ�Z7�������_Iݬ|�f�].m"X&�N�e��g��H�J�`S}7�!;�& �.Q��~a�Sȫu��z3=P��"�A���3\�|��"������ur9���t4ۻ�-"�m���|������}�G�Y��O��b�P2�<�cM���"́Ǫ<���n^� �A+v�y����&Z0貢���:6�`a5����G����~K�����Lo:��9�hG�k�5*�A�ˏ9R�a�)P4 ���$Ix.���z�y�TW��b��,v���4�+G�� ��r���4wZ�\N��U7c���Zxo�Y��Jq7�l_��Z��sh����[9ʫ�eVv�)�D#�3`�R�u|ǯEE�h���ɚ�Įà��g�NW���$���e��'@�e��	�AR�/�]�+�̂��-�/8>��l�Nw/*>(Iaw�󔛠�庾&��u�*�GbYܬFIj��z�ɖdG�GsJ?d��k"2p�Z�]��^�����'��՝�L�G7T��ȼ*����c�cb��3��۱�֭H����|���V�@�$TqlU����q�[�*�qˑ�\���q�o���Tc7� �!�������m�&����"`��m�#h�D?��?��+�;��S�3���=���/��bg8N!kL�z��v��'���B�oQ�����0����.�}s#?�Y�(�f@�~�)4E �HX��4	�'����Y-c|�j�98��N��\`~s\H�X��a�rO�V_V2��b���y��͆=��$�[ϝ�W{��oG	nV&��:�U��ٷH����j>�����b�e�`ևѕB2�a�;�&����,���,Jn�XH&�K������Cf�^�}֨l �D�b;�ԁ���Ikb��-�C�@~|�1`
)Bй���O/�����a���.2TsهϨ���G�f[�$��f�Z� =�V�����KB�dY���^�+\����-�\���K`�k�X@��	�5p����)��/~%Z[[v�c��\M9�3z5�� /v�G�!Po�=֌���=�Y8ڰ�/��p���_�A�}"�;�s�5�5�?�E�����'h�/a���L���w6PԈfG	�� �� ��
]����m��� �M�m�|88a����W/����5v���߯.>�`FI������#���e���X�Ά�,���XBR3������Dx����-Q���������z�P`���RŎq�eXA��+j�V��~�������u��,���-��3����D�	�:C�g;�$d��f�� �Í��H:~]���XAK�7���\��d�D�{_�u�.+�ǚ�����ڧ�`Z�i���nT��G�������B�}2�/�o�����p|���L �IS�>�ۙf�渌�F�;k��XR��s�|�Z[�Ke��j�6\�Ǚ��Q�ݳD�b�	:������-mf�iكu���%�*Rx�%�d�o�:�d�����v���)pS�Db���B<����!V�
3b�s� l7��,v�ʏ+�̵�y\��=8��y�!��br pzDkvY�����KA� $���QF��-�D������%�G ���Cq����X�������~���86�-b�1H[�"�J���Kj˦����M��/��W�q��"K�D�l>�O%�"�ǵr7�W�O�	��e�E8�E��<�z,�V \��;D�*w�����{s~����h���]!qP��|�U���RB���p\;_HA�`��+l�.��r��;�hA�+i1�"�ل���i����~zE�}�=^g�WtK�}*8Q}�T��C���1��r썽0{a ��P>j���p݂��zq4�����y�3a��0���E���$�;X�X�Jk��U����[B�����ķ�c�С[��
&&�`�Ct5�G���-��[�w�޵�ciY~�v&�K�*�?���) \i픔6K\pA!�A�;=�����L;��9���9{d���a�9w����W��lF$���<þ��6����~��p$��/���7~]��\xR(��5�rO�K��n/�3����ҹ�}]�Q\�OKAr�ʹ�S2�;B�(��_)��m�F��Y�]U��(�E�Y9N�r�( ?d a�.tz�^�IZmܸzO�F>s����P�<� ǿEr��:���q�׆[�w����a����"�;�o�43"3���;�[4��1���#n�.�l675g?��s����u=�SS!B�Ԗr�0	�=��^nhi��e��!j-��A�D�m��@mU���;]!���5ȵ~��6+nG���A��������j���Җ ���^�����͢5���4I��Z�����߅:��̡"�.��c.�������j��0�a�+�Ԩ�~�ӯ��}T*�i�U�]S� ���K�}���<!��~��.�%���N���1T⛺��0*�Y�N�N�֞���;��S�>�
��e7�����wLJ�,%<�xo�رJ��qi�uYyc���4D�tV�#ǜ�� ���/5�������/��Ҟ9�� m�z�VReԶ� Ep��9�0@!EZ:�x'C��O��Y���|NR��$����.
��/�q;"��<g�H�� �g7�FvVʠ{�Z�8#ݠHX�K0a���q�n�pH�cGi���TOW.Vr��'m-3&����0�\PX5b�n|�:�������Y������z�~���%3@�0�� ��`�#��#�����ެ��8�Oʗ�ât�^�/��2�}A���٤6�^�Gv f��Α��:��l;�˭��Bve�H*���AЂ��Pf[�!d�m���H����Q����8�Ux��N��-�����Ѡ�%(���u�*���0̚�١�)�`��5 ����N�j�O��=��+$��ڣ>@J�H.puFh�g�v�f��p�`�kK��F�H�I��i��.c[a|���n��W� ����O�������*+��L�^�-�]#4��i!� �åJ� ��FUa���j΃�_��y5k~Ɩc}J�G/=����f�n5f����떱�yR��2��^ة�~T��D�[��Eހ�vmm���=h����0��(�'��Tԃp��AD#n�]Cf��q=@-�1��u0�9C��'j/K�1˚�(�I 0�)I�ΔꛃTe�����~�F�Ѿ�%0�q42��R�_ �����R āRx��KS�	�v	<4�+�d2W��Z��X�͞���/m'� ��(�^���,.��Ѕ��$�l�W��q�{J+��cgg�����K�\�$a�8H�z�\N�sxL*�%�������nn��}Qv�ɔp���ԫ=��	:-K�A}�"��9eIfXX��V�}�����S����������@X�A�:�����$�*N\L����4�i"�a�$�</�ΰ������u7���Cù�[�R���P��C(���k(��g��%�Z�l>	r#HoE1�t��o��.G"�lxv����Z��M؋K�`����=9�F=���{�������~����E�SCgcxGs�R1/����:V'Ya40�^�W3����>�;1�4�[x~s�ډ}�Y�=��^�v﮳@��Θd��?o��Fq�����C�~;��M<��ǃ�tj�-��@�<̈́X�}��%�Ӯ�\S��}D��g�<�G�cU���*kUъq��r�Օ/�K�

��>�6�+��=��BN���s�>q%I}N�{Ձ�H<No*1�#`E�u����ڔ���� �D����"�VPE��<������MИ:\�bȠ�b-[1t��az/����W
����^��������?�5���/U��?�YW����z��L��s� z�\��g�w����T��:XN����q��d+���/Ģ���r�B���N?󫳌[E�VL��W��r�tIjP�qM*�?�qtW�ْZ"Q�?j	PIh�P	�^�=c�u���@0����oa�6�LD}���і�Y>ֶp�JC?:���79�g�y���A/8���j<��^�y���j0E����i��x�؛o7Yi���O������p�A�8R���5���j��[�3�V�k���Բ����B^�����盘M�vgN��}sG���|��4"�J&�%ʠ%ͳw�I�p���Gڸ�Je�a��$�ӥ6
w���r��s�m�g�
y�ac�˻v��Y\0>*q{ګ<	�P�/��|��,4&��k\!�K�a��Y�*�hâH�����(R�'l�)��:,��C	˖��J0�ś!LC��U��� m
�2����� {s�B�����^m%��	��~>��"����>�qV��W��i��2�G[����Z��"�<ّ�*s�;��s�YEV�)7�MF�OYX�ñ��$�G��	�ȟ��</Ի����eк��r�p�Ӟ_�+]�������B���}�@���R`�*ZU��WI�-!��#}��I}14��WA��O26Z�te��^}0j�d�w:����y�U�4�6���T�׽���L�����.�lW ���5F���("�ەq��^�O��Rd1˨��`��_�l	���uth�ky�FϜ|e�N�0�T�:>���y��'q�RK�"�uf���|��o���[G����g[���������e�(.�TK'	�ach"!�ˇ���q}�M���cX1�f��=��P/�=A	��]�J�]V*��b�D�A��zM���B
37��Pw\�@�m�7����Z�JS��cA��uEbT�T��j� $]B�����p��.v�z���F/������"I�@�Fq5��g�r=�f���f��>� �T��&���p.����T^���TZ2����1�C27���Ό_^{՛���2�����g"f1kV�9Th��ώ5�`�&B-LN"Z����������#�B>rIFM,9
}>�t7i�����5y>N*jZ���ᒴ�0��%DxqZɼ���Oѥx����'���Y�~�d�P�κ�2�F
p�s�#'����\���0�'��N�V�K:�]%�n��z��C��� D�[5����oC5�����ύp�p��蝅䵬!�j��*lY�Rz�1�{�K���c��%�O�����hk����&p�&t��"�w��z����z�N�s�Gνqm�~�#�ar�ǳ�ͳ:����� -�WP���Y�W$��mn�Y)��uS�-������V�Z�5<���3�5�ײ�\R
�| x�!��Oa���hJ����� �&ʄ�5� ��j:C���e��g݁�m�ذ���1����jI�
[�J�D��5.���\.|�t��L�T��h��?���aeb���wS�3s|>b�@���}x͹�L��D��ɪ@}���P�3$e래TbN��Uղ��E6�Op�8c]���l��B��?7�
�݋� ����E}�Z�W���k��۶�Yc�R��f���W�f�\AO���F�cZ�)��N_��Ank'NS���-`��i�R���GqC}3̜�ľ=��zmd�2��vh� �e�������T�gz=k��*{<� ���DOD����]����[���'�F;cQ���{�?�?���@V��y���{cM�
8�a���2��+m�
�#��L��Á���5)��'��L�b��{�>"M�����Of�)�E�	�v��f���l,l�d��YĿ;	��($9 =��SMR.ja9ؓ�r��,c12n#jLO��ϧ]�j��J���僰����i������õ��CS+&�ŀ��vg?%˛a�4Dy�c���L�����Ѭ�YOAhg���1�Z����IK��/�
��iTP����y.�H�@���:8��O������>}�.&� ��k��h�y��2�$�P4���y���{A��	³�Ax>6?{�P�E@���Z�� 7+��� r�����(9���c�=C
���?�_��Z���o�C�ED���+�pī"�9��^C��7V�G
���]Z�x��;��7	��c�5�4&`���W�c���OG�"m������Ma��QV�R�[1JKo/���96���')��G<}+�����V����e-Xt~R���1.�vij9��{�b����z�b4�ػ���X�'A���� �����J�E6�@c1�Q�z����5(\#�vu�d���i���(�^Y�TZ	���T��*k�R%�i���"�_Z	�}c3M���+��>�w� Y�ޣ�� ��oI�!�X�n�� ?�b<O�!:|Od�iC�ޡuU���B��T���*���:�c�N�g���k�H�q�{T̋!����)��F_a��ә*��|�gz�����^�AE�F�p�� ����m �K쩃���?6*�J����`TP�rfr>�"������%�|�9�H9��Y3r�n@�Dy��}w���b�g�5js��F��T�yR�]/'�$�^{�BP�R4�L�%V���z�C���a��f��`+={,!j��b�
�I2R����������׺��^�$QUٵ���θ�O1��
�N6��LA���|HAW�a �8�$��^�U0&;BGW�ݵ�u�L��`-��̼cڌn �mN4�$[z�B~l
��+`�Q3r(X���;~N<j�H���D�'��q�C���J�Z$�-�V�Q��=4�x�����m\�W���ѬoB��.��p�&�^�A����Ч�ni�G��O�Nµ�D{`�84X���;q ��E�]�U����fH�b�Q�A'��yx�ňb��~�j����J��,�"r�Nc�`ݞ�e�AvHhg���Fy�w-0��$]�ԗNU����#�m�7��g��In�E��l�=�#��';�_����\QZ�̠��%�dЦ}�B;���;��������P��aw�3�]��x�U�P=��F��Չ�XtT��$+���$V�&�Qy�z��^B��"j�dW]�H�)��s�����) ޖ.�o���=(����M��6��S;�G� =c�_���A\G�٘��|��� F�~�mN�I`T�|�P!��6:��� �B��Rߨ�q�w�U�CMOe�
�Ye������f�����{%/7��5I�xJа�n,_�$����ngu�e������;{q�!���������?�x���B�J���5p�2��?I�p��v�"%���E�����0Y'h�6���ǎ�LbW�{����][j4nw�:~�]��0cY����2��Z}�T�r���1��4�&�qJю��ۭ��}:�(
:��?��T��tk�p�Z�*��-S�)��%�6�d];�U
���Rgx�Np�@��U��#``�1�K#���i�M��خ4���Kjh=x������7�ei��K;],�5V6�0&������߸��JӀ�c5Dф�	���=�p&k�<���
sl����q�چ `�J�xB�!E�Z%<Un֍�����2�拇�̠��ɆVŲ���	�a(����(��d�~�9B�嘗c�޺s��W�iJ�>���/�<�AAR���U�6,_ kzL�@��e�+���u>k�����s��W<a��<)�����w.n����i��'�S+<����޺qm�����@�����1�T�G��`�W�r����q�|��RtN,'�H����[5��{M^<�( �I+A�s`s��2J1��t�_z�M�مM���6��{>�W��bM%3��-t�o��Tҽ8������C���\l2�����6k��j:Æy�K�~{�l��M?m;��.8a+&4��W�����t�:��ǟ��CW�i�V4%<�h����-d�/�ځީCÔ�Ӧӆ�P�+,!�~�x	0�D��,I$��?1�������kÞ�CنNs���ߗA�f�o�F�Oo��Uk?�4g����6ʸ��*�)�<:T���">	�s �5��p��^� ��7��\����q�����1�����&�B�o>�D��7��!�%s~-��|Mýؕ��'o㠺�@{M��P���:��p$���=�-���V��� /iM���p��۰$�2Q�ЖI��I�!��S��L�8��(z�����-ߞ�*�m�����!�����i�&��ǁͲ^����Yxy]2ߥ���n��b��*�z���&��@W\�N��Œ�@�_YQ5�b3\R!�s@�iP��R;A�����ڦB8��Ϣ�X��Vm?��/�Lݚ����GW�	��%T�P��:��tX��IJ��w��g@���B�����똳�	�ʧ��s�FN3�\F��wG\�v��b�N�1+�D�;���@�!��E�];"}T 2�s�A��ZJ�wH^�����cA�k���������B䉃3�#��_�O~��DG�}Ռi�͢i2t��<�9W�+>V*�\�!��$�y��
�~}���~�s}�44���(��v>}�ʰ��2�"QT.��`{��U�o�5��Ln��ϭYIVx�3DS�9w-G YB�3��C5�e��է����FG_^�y�K9x���?KF�-7�D`��{�[bd�#u)_#��m[<{�$�����(�����=�=	�Lµ�.�K�E����d���Ec�����F �ד���~�����(�h�8�B��8:=�f�/�ㅨJ����. ,�܉S��u͹b�
l��:ӆR����'���sԍ�\��;y}�G�����K56��q%4r��' ���ɒjF�F��b?r�������8qo���kJ�l�b����%~7��J��w 
�4�A>��O��^��D�[C��C��
���F���6E�(N0(���Ѭ�k����kv�b��iՌ?|r$ga�gz�S�Z�NgM�I$Q�xW�7�e�c��5J�h�C\]���>�ɋ����7��n�`�j����"
~V�<��ʋ1%P ��k�b�N�i.{n@5���/�؛�C:J���M���QH�����PO�1P�r@ڤ�ۓq]����ȯ�ފ��e�_�1�w��t>P��'���t�r|[ >��3�=���|,v]+��!ceq��q�Y��u��.s�r�r��4�JKc�T������7�-"�B�����#�N����qES��n�����W�����R北0�W
0�q�i��u�3y2gf<Q]4G�
,2�y�F
�@�/�VX�GQc���iD�A���O��D��;se��y���3W-O�s@���� x��:�z�ug�kJ���Co�#p�UG������~��b��m�~%C���"���SlYe���N*aW� �q�'�<�ChN���g�J&oѓ�ի�~�⧥���Ox�V^I��n�nUG�W���Mdo�5���8���R��mQd�|3����Zr�������!�%q�>��Z󗼏Y�~�gYkNZg(����G�T'����;�b	�����7G	�Q(�5ْ���"�}��N�w0Z)��ʿ�3> �����h
������P	��>x-��P�;�"�_W�g�	Oz9������$e�o�o�`Ϭ�ڜ�%��)��fJj�z��_�kx ����`��F�,�Z�*�L0^�H^Y�02:/[^K�Y]|�TPK�cjR!V�כ��$|2��ds��-+�E��^�5^J�/�KҠ�a�����Sd���D}(��P�P�uZsM�H�IE��[�hjSPs�����z�@*�/�VD���I'��rL��ĕ
�q�w��B3�^��Y�W�f��;���>kRM���QL@�����{��3~�B�X���RGA�#�lثx�c�,�Ͼ�И�pμ��]����W|p� �����q7�gh+�y_Vm��]���w�l
ڄwf�N/�ls1��C��<�2���7�@�'<��f�؜+*e���3�	����A�L�6���=�bW�T5rzy�������YO,[6B[�'�H9��}Ӱy]B�J& �עw��Ĥ^�h���,X��O#���u[����qeGd��r��B� ��P��֨G���*!&����R��2�6oHK�+Y�"{roȋ�ՌU y����=o�y�xA�������.��j�B�y�����a�K�vʍb�� b���גe�u������˳��F�ֶ|�$�<�� �c�z��H��QT�nկ%�Zs%��l�sK~�9��q�Zd�L/��9�X΄�jY���!O��G��R.M�?b&���ې���(�L�������<�>5(��s30J���ֺDB"�`7N�� eX�ތ^ط�qs���O ��5�k,�h���i[8X�.8{Y�e*K���ѐ@0��
�(������LJ�Z�ln���hó��D>Kwǡ83�x䡏+���I���5����.��c"7�B�aܼ������[� |�����1ӫa�5�������&~��C���8)�A)�䰞�c�M�J��X*Q�Wm��8��u+FD��d���6�h��p���F��>���,&~e!r�r7"��ӹ�P�/�@b}dN���T�q��$��}$
���|���%���	�(����yh�S�K"J�\�J#3�FWS�F�&�Bhq�6���4���mz4��:dPS%b�+[Q�M5h�v1�:C#�=g0m�ki W�Fx���U
L_~،�/���Z�K����=�E�ɘ�G���+Q v���u��cb"�p/	�����"/Џ�|�n ^�9W�DI�Ϙ�^	ňk�	V���ݜm?j��,���c;un���#:�`W�#���\��a����+����1���z��MX�τiò����m+��M�3	�����S���� i�����d0�����=߮GY���;��P@1��_����{ IV�q��ł5�l��+TW�'�<�Ϋ�ȨԼlnt�e���2�B�,���)Z���O,A�,|����1�U/Ge��l݊����-j| i��o�l���tywz7ƽ�������\�;P*9�Z�8���~�n���lן5�S��A{'�m�� �W���$0��Ud�l�i��0ګ�ϒ�?��F+>��.H�\�t:��5+���2�(ߞ*��2��%f�5S�ǎ4_��G��*r�TPz$�U�2��3�������}�B/����k����FB��|���/؁	�t��yh;Im'F�q��ʠi88X|��m���*#��tP�n�ϋ�N��|��)��NU���q8t��4;�q^���d{i��i
'D��P���[�]I�߫��r�('d�3��mh��,��c��"WS�%�3c����gV�7��r��ҰVP5�+���zܶ�^'4p,��du�p��|�����JQ���Z6O`��ܜ�_��Ps�u�B������$�&�n����,��sM;���Ϙ
ߕJ%���L�rH�~i�w���q�p���T�4��j��ID�hΑ��6&\���jR�؂�����N�de����5K�@�:ҿMh�~�o�%qO�#�H8��=�qox��Xz�x� ���ڧ���S��:��X�stG��C��y��@I�D@�4�(Qh��|��}ͱ%L*�/�B���-C�2$�ډu�5��=`q־���k\��oQ�������B#(���fy���/�ҹ%�ԕ7�E�t�]��r�
Þ\{+�_�о�\>��C��rw�ۛ������R�M�?+[���gt����jNp��t���-���r�\�[:[�}�����L��q���D�ʡĨ�ӹD$��ߓ׫R�X�u$�B됿�:BLXe�U��i��%Ю��/��y�8�&f�|ڪ�<MSg/~B��ZF��!�7)�#���޼PO�	_G@>&�*3�
[��:ᵓ�{>�$1��Y� �F��V���~ؖ���N+bLE��ls���j2_��1���ky�틒	�i/@�G�A�վ��(��5o�!��k�>��-�F/ǨB��VHh���`$�5�rdh���P�@��L���k�;{fW��q�*��*�0����\`<��n}���:ɡE��p�������������/�,C�Wz)�h��5���oj�a�o~��+���4���M��(����
�+?�3��j���X�6N���P��:�_��z��>:��qjs���{޷9�B��ϳeA������k�驘�2=l��$�[���?�RI��*xb��h�e����eye_Dg��){F#�Z{�)�����7��T�%�.*ڋ8��\��N�W֣m�rr�׽���$�x���F](���H;��T9%�N���V&��ub|Bf%�?�W��0�Z)K��t�5x۽�vՆmծ�B�Z�I�~��O1z2�*d�w�j��M_�k�,&i�VY\��L������a�ޕ؊�=V�V(q�Ir^�am��҈*?^t��GI{g�'����%����q��5�{�nK)�����!�T��kE_�F|�ɩI���vg*�?͢� *iS�����5b�R�<2�R�ㅇ�M���C��O1��q��z���,)!��䨿�銥�eyr�;��#�z"{_�]�Y��/;�N��s�IHKd#$R}��������L�@�/�����ێ���(��.�%+���};.g\�@���5�9f�;�\��7{�lK��BC�!�{ڐ�|LF/��V���U%�Ѩ0�!6���l�.Mb݋OTG����|_��ai�p5�f��V�fNu�AAM�9�#�+�Y�՚�?'�}0I%g!����a�v]5L^r��歓?�y�:�%wt���d�r�;�������n��<��Up��g}m1`S-w����U~sױ���e��0JX��eŰ"3B���з�L��o}絃U�9�X�S����b蚄Db��� ���#Γ��izz�Q���D��-l�U��P�C�Y�`XИ�q���]��8�D�V�k�C���2����s���}Z恐�2w�0�R`(a�4��S��w_;[�Q�������� a$-1��L���h7�0tPﾴ��D�ь���P���>��vOY���&U��[��KN��]���31.ؚ�FhDfԋ��'B�t�&v��ͪ>��{�< ,юN��y��p���@#��iթ�ȹ̅��km����;��խ�����%��5q���{�'ǣA��!�r7�iS�%�?�kY*�7�]7��'���ɱ��+��f�@�l~Z�b)a��,9�X[(��1�=E��`�ߵ�k�4�����t�.�G�)��
� ���l>�V�/J�^Mo��f�\�[(WQL3v���ϊM�gQ����)?*d�iv\�އ��M�Y�V%H4�YHڒ�� ��3z�f����{v�p�li��>{	ӪF�����>���&��<J<8p=����j2h��ο���/R�l�_bi��8+D��^&�ф@�����=Bȵ�>�JbT����H��7�œA�d�#�:Ȝhg��ؐ�ϫ�q�;_��V	Ǟ�XaQ�����$��X�SL7�(���fE�龬���S�FG m���F���������3������ޮ��+�^g�!�G�©4���7�s�q��r�]�c�����c�P#
�;Y$!/���_�7Ԏ9����~�M���X�����)�X�º���R����͊�K:������͡��
S /ښ�]a�oC��s�'��4`�D+�ɱ�`��w-d��?�������xl$>�	��h���JA� I��+�em�}����`P��s��s|�0�]h*VA�b�
\k��`�*P�z`"����K�qa6�������zi�⩷���� �����'��5o1��/�ž&u��Em]�6H-����xcR3������/؋�bw>�Q��o�O
'�8��9��}�	t�AbDX�pE=���+"����L&箣��4��ǐ|��?�Wᚪ�Q�?�`�Ђ�w�Ay�a�	�3�SDۃ�������Í��Oz�%�܉�C�6��HǊ���VW�nn��oJT�5�g�A��6�W��Zd	��B��]P�����G|@�����%U�2	m!���~�O(��O�=���L�h��|da�YԔ��m@�b,I:+` �gEB�L��#S�6LO%~��,�e��K�]��p�P�8��A���4V��ԃ�-Z�
��Ճ	���RN ��9L����������x(d��a��lm�O��'ET�0�w���[gn�s�k�<�J7�Q|�$,]��9	Q���vؚ�=��(��$��|�����*����mI˚�(�E����M:"�}�d�"=����oL�4�}�rp�~3r���S�B-��Z]�f��W�j �d��!�[���f��_�o	c����\T�a���Xa��C;�#��Ȓ������(c��i����w��j}9�u5Pk�_�x;��h��ҁZ�(��61R~��O�I����I�S "�k($��J��
d�[^�M=��� �?���:l���4jE|����s�:��������Ξ�wB�?!TDqا�$_/[{�8v�[*��W�IB�m3��dϏ�!>*�/��7��f�bG]�oA��/͠-
��G��iX�A�h���3���!��[��������䩨��'\"���%��n��_Tt!�kmL=}+�M�1��;�xGW�6㙠�Ɨs�6�uQ��d�Z��'P�`��qҡ.`'���p����a��vk�`����C�^��>���QTz�dI��>2����g;�eV�-}Z� �Y5�y�,�������h[�7�hY���O�,�D!�����B��7�U��n��.0(�!��B�6�mv�-+t\Y+�Ȥ{���A���� Yl�Y���NJ��e~��Ж����ӄI �����O{`��;#eYwK�a����^:"�O+���d�T��WV��jf&���ŨT�6�ld�'+M��4u��͗����`p9�J�\G�A�p�����4���A���,�k`O�$B@�tIA�A'�����BЇ��a��>�w+�i�ɏH��z��{!�}sO�*e���ۤ����&-(2�8΋/�Ĵ��4����a6�U󳛿O팧L2� �69W���K�n����c�rl�dM�q]��)_�
G��{p��*��4�:o
O~��A��p��K	Ý�*8�;!�.�|��5�a�m��Y�d��0�V��n��rS�z�2�ZBF�K��Ji���Ny�W.X}x����^ 5�wY���!'�?O�PѮ�!�U�4��ԑujp6ۯC��m[n:'.ĕtmr��[�Y�����+�l�����M/[]'WDἌ�b��NEKgKSK�,���;7���7O"�z��n2�È4�Q^��D��~<��n�{��:ID�]K��yZj���]a����g�\F%�H���D>��N���b�:�Kh�u,WrZ�!b����Q_��)S2M�H�N�X\��(���!	E���^?I���h�HpH-\�b,v{��"\l��4���u=�u��`�j��՚@�y����q���,��/̌J�GY�uaWs�k���_��5��_���+�D�䖔D��:��Ti�H�OL�|-:����u@U�X�+�p_��ь(TkxE�=�G=�����H%����5�\M���A��"�Pn�-�nP�6���jΖ	f�3M�5�66�I�)r^~���<4�#�t�mV��>��~�*������쪛��AHT@wg�]<:��Oف9�*+�����9�J:�]Ζk��r0OFѯe/��0��&��kN�i,�x�VBMz>�g��>�,'�Aϼ��Х2�� �"��� �u �
7�Yzx��8���	�}̵��?�:S9?¦�e�����ߪhK�M���.!�����J��Z�����@>�qR09�0ݘ�*�#�+C�8m����G��P��� T3϶���'����j<�r���䈼����&~��[�3U�J��Ͻ�8��}����4�%AMv#�j19F�)O���/���[F���_y���� ���U)F́���
�tIOJ�{ߚ����T�b�[Ј�?���
X9p�b��xC���p5�'s��e�ZH_��͒�:�L���[�Q���8�I�IJIO`�sU!���\$)��D�\)�u�
��+�n���e���~��� ���Mew��'��|�.�|{�l^
6�s��(�� 0e����<�[�ج1��
��S��1�y�i�I�v�L`�g��m��Μ0��D{t0�8MB�U!qj��b�y^�b>���o��eNW��%%� ���U��"=Ԙf�K$7�e^��y_ K�f*C��]�@��nطX��;�w��ͨ���-�����NvnM�͗}���%k@u;�bJ�T��o�#����@����*���	��̦X~�Qs7�е`-����ͽ�l��v�ԉ���w�@��Ru��o�SƮ�y���ېQ]��v��s�暓_���g����S�ަ��kf��
h�}��o�"QWl]�RR޷��4U�w�@�ҍK�����An��?�j��>n�lU6�hN��{~������f�K�]љzp����iK��ڵ��gB�+����=���X&��AYy��e�nk,�Pm���p!2#7&)q ��G;b��"���x^A��#��M���="T<�h���:����O�I��!�Y?�T-tC5���:�H\!�3 �ʷ������%��3��������� ��4_�xP˭�!V��[��M7Dޠ�ى7g6��YJ�6�	�Tųa�"��Z�Qs7X��Ѯ�Kpd;o_n'4I����73n�ː�Dߙ�#/kp�����Kʛg�[v� ~]v��BFD�1�I�����������l�DQ�?:�iƈl��-ǘ��e*J�X6�*ho	�q��nz���T�f=��<��ΰ����!�/��P^o�v7�k�Q�/%�5�Zio(/遒�'��6���jT�<*����4\����"V��9�w�VgQO/����"�/���E�ˣ�47u9�S9��Q�o�M�->�#rP�SX.Xw@�T ��R���F�؋��z4o� :�.��o&/��-�n��<_�� --JKs:�$��D�E��������w��!Y��@�jF��U
� m��|��O1����X4@3�V��u��Q��]���֙��5���{�_���$t�@5�s|���i�qz
�=�Kq�]��y��|�YG���ʓ�w�YJ坖5�Ū��o�[������q���~܄�\}�'�r���6Rqy	 X�������9.���P9�þ]��N�"��}.(+�?A0�sw�a6ϕpo���\�+5��b�,p�J����68]Վ�]��_���z���5�r�'єY�~^��@**��r� �Sp��;�	e	�C��@pkj~��w��.0=��i���V�k_)ɺ�B�BG(/��Ӎf��HͨH��o��D�4���Y �ÀPJa��m���A�9o$V����ۨ�/�F�Le���[7���7��W�!�K��D���	�H� �!�I<��U<�2��X���KT���`�%f��¡��W�O��)�l�n�]���(�X=6�wc�'�g���^����e���J��Z�c�D
�T��J�_TW��� k�� W��hؙ9C�&��:�]R����9�Q����*k�v�8��_�A�lڅ�N��G3���+��!��b�
Q�2{䰄��m��B9j�,.����U P�D��H�z��l�w��%D�Iٌ@�6�ZRG��b�q�v���J������U8Ú�H���z�
�3Ԥ틸`��x�2���
�]^w�ؓRd�î܉������#?��?M`F����Ǎ��'o���d�G�b��z�=�n��XA�[Fc�TMP�LgSk]/c�d�O$�T��> �:^m��(��R�[)Z��� ���e���~x7�fxu�UC,�%�I�MG�k	Y�6	��o��N�P�[�E�%�ӏxy^TP��{�ȚPj��R�&�*#0ψ�c�s3�_�fR���%�����мQ(���X��o���ɗ�)�����!�Z�>Չ���W�%D�X�w��z��ђ3�vK����ʎ�5��}�;�E[�Dbt:��S��lc+��ĎB��Bv�uf"{Jb��H2A��9)� /+�Tn�_�)t1)Vo�R^dv��EJI <��/4� ��ӱ/U�@��1�� �	�,Ă(��?:�z�Q�t6�ѕ	��e&�����$����9��%�mضG��j,���z6k�R�<a���	�B�*���It@*mJu;����C�@���ٯ���3�:}b��޾t��^�����/e"r��Ɨ�G(دSe�+p�EzW�A�RrH��e����' N�-ß� �����'�@:�Fx�j	��d�����B�j��ۗT!�iV-�,�}�V3隌{֡��<���k�$��%��Ww.�9E�ř�B��Q����#�ZvW��E�LW���W�a�h�D6y�z+n��S�ྶt�������g�b������L؈�� xgvK������YX<� �,̬���	9�r�m��cd�Z�3�Q}T��g�x��������E�R.�w��R5Z��J���#�������Z��l/��Y�k�H
M�G��h��L+��^bc� �D�ڳ�	-��6U-�,��X�V��l?��N1�J
w:�N�h�:�)\U6RQ0�o`�1p%�ÅA�}�rм��ǳ�^��V9�ͺ0���O��{[X�"� �&SGԲ��7)u��=�]j�����E���D����b"| ʯ�����p��y�P��p� '@g7�l���>3.�g09���K��h�]
B���4�.#�ܩX􄳉��ps�/��ʜw�'��;�j燜��iu3b��@�
�T7����S������/�����*��PF�Ij�|��|Yߊ5Y00��t�(8V�Ł�*h�hӶ�vX�
�W颕t��P/w��.0kz����Kg�&���4)L|[ɿ�V���������[`�P�8�"2�+,8����.����P��˒A��%X��ݱ�\�e���yP�G�T4���
^}�h�e-Ӫ;���`��;�P�a۾�3M��~VC�0b�f�&��q� �9�i�� ��q?�=!���^�.�8K�[v�T��T�����I�k�j�l?F �1@6{����.����V��oKW;�O)��H�.R�i��{�2e�a�|�ƺ�{?b{������	������>)\��*�|�|2g�Z���M��D��+Ѥ���9��*��)��!2<�ޭ/(k�w��0
�Rl���95��l��0��|�ܿwYM����,�:*�FρzlY�����U��6pa�4��E2Dx����S6ɮ�2?�n\��W�o_��+��n¸������3���%��r�V����w��,D�3��`cbԷ)5�)#d���k�H�q�?��.������T, n�;�������~6��&\]����C�h�A�
����j2�x��y�@⠎��#�$��������P2�����vǌY5�AM�l���7S��h$��G�(6XM�N2�x����?�oS]�(�c��3��m8tp��n<�A���4%w���C����Dהr�z%��r铼���e*h��S��&g:��9�)���=7.���Q���{�a}eq�@��u��>։ ��c�Y�pcK,��#�wg����Bqg�_���]�5�ad��{���^c�		��e-�R��=R;��^Q�x��-i�D������`�0S�u�Xt?}���i ��+�a�]��|�'��I	餰�)�A��(�3�&��e�XJ���p�pzY�z����ܟLqN��Q'��qq�I�L�ԐFW k/�P�������I������֏b�C���Zf3Jre���F�9\�0�����5x�,������'���g�ֽvNG�/IqwG�������~����K"������4���������)<.{+���-��1>�Vb�h�� ��#|����s�W@�Ϛ�� h>c��d
$kT�=�K+�b�-`?��BA�|��ĥ��\�'�Xu��·,(S��K�[v�mGp���D+���^���rV£8���&\c\$�5�Y��UXZ����A�b�������	:�F���$������n�5�\�@m���xm&��$��D/��	��z��;Q]�;����
���s�a0���PV��N/�ѿ� 
�F�u7M�U&��</o��kw��-�MB�S�����*(z$@#����3�g7���&aRZ�6B��7���&�t���R�%}�ȇ��V�w�7�&CwD�w1����MgkG5Ҍ��PO�7�����?!#��s��1��b�P�C�I�M�U(뙚���M�^�]9���c����+ȿ�2g;o�fS}TbÃ�7T�AU#o��:�G��Kɐ�:�ji�nSEOg<,.�z+�zEZVA��1gA��d
P�v�l�8v*�C�L�����@��o#x6~��jIx�$8��3����jH/c%�%`wI��gЋ�v���P��K�[�)�i�*�����saN�r�|��V�����L��;��׼-�N�����mT_-oy�9ħ�N��<����p>�}u��-�j��h�V�|��r��س/)�8��w��W������&�wh@�n�_��<��6u�Ǐv2�P8�Q�B������'�[ϜsS�"szE~�^��B�6>/�-�w��m���.m��n�.|*]��K� ���" V[�p�2ߒ�L�/��
��$� �|�;��3��'/-�cU��3XQ�w"���d�(��~��iG������*���i٪�JSt�<����XMR��0Q����7�����ֳ�s�To
;a����j[�����S�s�.Ц7�T��CLK�t��X�Sn�&I,��F-`\(�"��Q-��w؉f�/x�s��ס�ӭ�W�D��DPe�>q���eM�]����P�y�:7w�:���Cz���I� ��`U�PN�|�:F��aI^�'a;v<�#R�`���5A���CX/�
*�^�Z�Ɂ(>��50���{��㨮�Bj�K���r�ͨUtj�A��"�
�T)��t,ө#���՘N,܋/��&��%��5�W���r�#=��(!`�2�O�郮5x77��H0Pޢ���%��.?qD��I9OGF� �T�#�����5k$Y����2ԁ{0L����##��h��^tE���r�T�9�!���y�"/ױ�0����F%��PKpʁ�C��'��I'��S�1l( ���<;h�
C_Iv	Ļѩ���]��@��o���G;U��\�.���>����|�Ӷ�:�ۜ��q �E�c��q���
E��3˜�Q�����R�w`Of���")�C ʄk���SלaX^��%@;6븎]��)�n�_K�4F�D��&&����x�F�=\s��	2on�R�ȔF��F?�C�[ �03H��C��k��c�F�'��ܖ�ҧѹ|�}��<v,
�د0Z�Q?��
n���yD�єJ���~7��T�(�/��aKk�����Y9ա:y���x ������I��� ��Z���'S7��<A��Qr:�����-|�]����0ϗ�ݖ�D��Z*ѴҔ���#�g�=�� G�ݏ9����/��/H�Uʪ���"w�N�O���S�FL��cތ��5mѬ�ώm��N/)�/{rο"&���#�mVG�����7�R����9?�dJE��w�d��̕HY$Օ/�b�9��'�f�|��a�w�<�غ6n��'�(�����Mb#�F���r��4Es�*km,4y��Z�Q�<UeM�Q���Y��WT��#�*�=/��r�3Fe<���'���ض�z-�������q����ˍ�@:6��I:�6ۄ|����[�i]_zwy���P�z4�O����u1�M+�꥝�6�&'n�_�ogP�s�o7�,��K-��?�!&d��US��M�b���C�]Em�6 �f|���9Y!ď���{�����x���$��h3w^�-��6rl���������2i��]���ؠ��������O�`��?��ϻ�z�Adw��+�-(oˌ7�(�Ig�ʓ�H��'�����Ml�vN�<u=:����
���KҌ�#�",>�����d=oQ�dt�����⟃�lX����3��l��v^j1�ɥ-V�{����Qֽ<s�o�����[���X��i`��f��s��c�S�A��91�zz�4ҧ�|��9X)~�jv�Wa���a*�Q&%b͒#I}D��vh�-)(�y�K�c���'>���KT���P�����$GFо���a��
�鰥�+���ȁJ�zr��ЩG�Ì��cI�v��g�ތ��~�H%_��	w�����O_��s��iO��n3:����;b��ۍ�ڧ�>���d�Í�Yd�B{��Ȟ^W���&����s �:¦v��Y���>{��s�'>B3h�UI�r;?]��^'���	�h�o�j����Q�oN��ؽHG�({�~�Db>f�=���S|ڄ��ѽ�~W�x�y��K���U�[���k��Ŀtv���B��=!`���\���P�ۼ&&P}R=�G�TĔ�L)ײZ��W+|�L�)">w���2�xƦ�D���P[��Ӡٔ���vK��g_��7�J��gJ ��y���;��`Y�o	_�񲎊!A���k�>$ti����1K���0���x�9g��i�1�
�6� -$0B�KB��TFH��� ����h��S�ؖ|�U��r���ߛ,ES�BWg8���g0q��6�>%��k!q�=�����G��Ծ��I����u~�+i�̀8�<1�3/l��p�@^�ǢsAL���6���N�:]�@���ki�@Y�X�F  ��*�������+x���|�d#�D5紞�B��s �覡��Z�v��R�1n��L2�z�9�p]R�������S�ԣ�4�P�{%���DV�M�x�עV�SV۱AU�/K|��r������8\M�����<��z�\<�r!d��o��˸���k�[�8�@S|F|�s^�{P�t�Z�x���?�V�`4���0��N�F%AHnʡ�����Ʃ`�������y������ T�8�ց���K��q����ƣ���ʀU�L$
�c�#���T�������"�� �]�r2ܺY�?���-�8\���}|:!��I<�ʈop�dZ�sCX�5L�$�C����C�_9�`�]b��.��S���Y�o�30!� f�D�5���P��` @�Y�7\�3��/�g�HddA�x�y-���*�U���O��
oX�
��B(�fj�D}=�c�R�/�[�1NC#>9n�Kx�w#��.�lɘ�;�N6����u\C�E¸v��,���$G�8x��0�sC��:=΀�SG���:I
����x]�uW�7CS��^\�I�C_���	!k�T@5�	�� ��B�eC���&�*���UHuG�qr���[N..�JT�MxK��r�+b�NhA��4��]��G!�"4�,C��C�pL�tL���~2y���)�'���e�O�d�8h(e�	$rG+\`o���J��3��I|�P�1ڶc������.�򉜟c��r����	����1���F��B�p==����RE"|�M(��d۰=���V��!#�a���0H�>|�-^m%�s
�ߘ��U�_�Z�)�+���gr������F#�21w����_�Hb.��h�BD~64���J��1i�+�l�ɓ̗947M�(κ9;�P����	�kO�v{��6��^�}�Ngr'|��[)�`��k��i6���pt�|�L"�+�
F�e�u2�+9rd�G�z�K6���Ht>��"8nu{<���ʀ�ø{���5�����&�U+W�17����_v<l>7�R�� �����2?�(�.�9����.Y�RX3Iv���Q����J�V�s�-��f>��)��	�.6]Z�3֬AEl��L>8[�5Q}{�dy1{�p�eʹ('݊g�=�m[�`�,XRO���O��9��Wy�����6	� ��Z�$w*�^���V��k*w"�k,Wն����>4�qr��j_�C�%� X�}{�mj7yp��ǣ<da 2�pk�-�P��$ %&�����,�ƚ��r�<�|�PA�OgL�o���`2���ɩ�����1�]�h�釕��T�2��C./�޿nK�Q�D��� F2�j�����L����o��}� �A�X������ΩR3t1`1B�����4��$r�+��!��)e���7��+�l齫
c�������Sxb��":l�������s�����Ti� zu���YèK�_X�}
�����$�zwﯻ���4�7]ݝ6��1 ��>�f�yw�?��:��ր�@���=�ø�*f��/��/�N��u��!XɊ^f^�q�Pe�ޜ}�_��#×В哽�Ib�o:�����\^���<�}녍Y��_���I:���m�L�ׂ��J�0�c��5�b^F��_�UR�1�	7�։'4������G�#�iv��)����N󄞍Ϛ>����g�T�t�[�J�ۮ�����A��]�L>�@�Οq'����(>�F�q�'���NQ��d�<��^��H��#"z@	c'%��d��@��kG:��"�Y�ưm�7�e��ޗ@�}�!C�.jh��1�X�4�@;��<������O�F���ij/�n� ��F���l5��AC��x(L�@e6���8̈��=d�tT�`�#�.��2Sl76���DfLACЂ� 
B�@�ԟ�?B6��t!$�:TѰz5��"��0�}B�e�i�u�Z[cP���0�oo���׭�p��n�󑁢#��CZ9���!!'o�)I���S�R\9�������FJ���o?j&��h��'���� j)��GQ_{mH��#��Y�:���פ)�e���Yw�m��)��^I՚Y��ҟs��"��XN��7x-�{��	1	Wu�~+�4ন �ُ\����z)0C�� �.\�n"�+�K��?�5�$X�O�4�gx�o�o������*�车�Hms�T[tt����_����@c��H�^��u��6F��qn�)6�>�k#��9��̹�v�m���S�E���4��Ǌ1�꤄T��Z���!R���~ʦK��wm;n'ՙj�j��L\�v'H��i��+���^Q�����l%S���q��ع������s�ս���s����آ�\P��`�G#�q.[���O,3~\��Hr���S�ɷ�v�W���g>��?4�N,��s������ƥ���$�	��P�X�Ө�5Ŋ@e���G�|y�эI��uI�� �p6�U�����*��bf��@]X8u���o�]�8�;��٦*�R�d���
"L��sO�����hQ58���#�����v��Â��H��VL�Xq:L L���K���ns�⭓�(_=�xy+�"1��e,z$C�T��	��C�i���F�bd�#�_���V*�ڢ�fo�툶���
���h����3ʽ8|,�ŋ�ʿ���t�$��jz�e�ܫ��PN}f�� 0|)��?�޿sE�{�	���'�(y�����W�/�k����yE;��I"����6�ʀ!�� j÷&�:m�ؚ�Ŕ��)�^���.�|��)����4/z77դ%��Q�"��)�w�t)1ŝ�Z�m��r�����"Z����6ؚ,b����ob�;`��:�]t#RUWV�j�C���>��f��d#��Z��J�d<�)�[�l�P-�7�[f����{�z �u�E��f���S�m�^eX��D�j���L�U��Ѧ)�P��n\A�rU�y�97�C���n��.��ul	X�/�H4�l��Pvof���Lӻ�P�x�I.w?\tz��:�4�q�Xj6iF2&���#[�H�o���'����3�� ��>��|�;/��w��o�uZms�&�^�.膞�����t�qpJw��_>~2�#D-O-K�B���#���%5����0+O���_h�9I8*~�^͘Q����1�;m���Wt3`�����_a=J���1�]8R�ӎ�R�-�e VO�>�Y^��O.�s;�`��ce�$��8���?�����\����;OV�/����x�ݴ3�Ԁ8�3u��� 4��Ѹ����2H}�XHX]����)�"��/ӿc�ǔC7-�~=	�WɉUHOh�$��jsj���h-�e���~������>Z,j�~�S���m�/m�1�����$�UC�/���k_�O���+I�&ҁ��v�^�=�C�!U��'D`G�JZ-	h��v4�GG��e)?M��o�b�^�g�������Efc�R����I���<��(;՚�F�eQ���r2Đ�����ٔ|A�R�K�U���N��2�W�Q6�M/�I>���!.��B�C�<����~3����k���VwLyFҧy�-)w:LT<�n �3
%NI����6yC�43<	�����c�W�oB^Gf��T�
�m��Z��e=w�)3���J����i9d��G�17Ks������j+��<��T���{ۘ���Tt9	b�5���!c�<��4k�	DJ_IJ~�r[�p�?��ۤD4L���l��Y����j�)�OY��QZ�8&1�|a@���݃$<�#2�8�J���z��lr���9f"�0
rͨ&�Nռ�c�A�����s9T��ּ8�B7(�{l��L*�Vi�N����;&��n�����圜BAnde�&N��CT�%�h������09Q�*?�Z��h#�0�W��+�Qd:�a�;!y=u�E�f����O�LBR�^=X�Ǘ�b��m�R�yJ�ěГ��t�tq��|��H`���������${7���Е��X���p�%qT�9���L�\�(rO����sru�K�����8�M�x��#	�J~|{qM��#����1�~I �Hd����RH ����Y�!�!����{��H9Dx�W��T�'���ǌ�b_�����^a���R?oB[R3�n�.�r�]>m��)��r:/�9g��G�F���.�!��R����֔���q�q�,�	�A�#w��k�k�nB��W����q]J.�;�l�qr�`_�)X�-;{�!�/ϗ=�#|z!qG��f��3O���3#"�v�\u�ޗ�}N rG{�i��Yo�W�S��9���t�̄���Q�����A/ʛ�\】w��%����c�a1�v,�'?��Bk���+�-�A�< W 2�� U������	��)&�O�/���Q[��WB��\�(�ݳ;��~��:�3�;�Ȇ�7������j�2�Y��©5����o�:�����A��ʞ��� 8a#&�&A�k�`��<ݞ���@c�W߼���	@���_���,<�qc�O�v$�PH�|���A	����!���ǂ���T��.�Qh��u��9a��'��g<�����X��Θ�y|@��#�cmFDu�_��Ӌw&J����S�Lx:��>k�Z@��X)@T�2��xy�?�i2�HSI�)M�.�Y��`2m�G�rw4�o��.j�����ni���~�;��1� ����ko`"��BB�'X꫊�+W�ǖ��A�7��,v�koWs�(yQ�ff�4�V�}i��"��0��9�����2=3��{�@���QSE_s��{�"�P����ɟ��C4a/� \���	�U�v�Z�^�l���8?�
���ǅq��P���m/� ��n��i��CP.
�rW1#�����\�.\�!�܆��Ց{Ԟć�|�������$ľ�QJ~#S48m��;�� ��16�)k�:�b�f�1e�&��P(�*�~��E!�(��r�Du/��K��e�Jݓ@��*A����ѳA�3����8bl
����V����ǖ��nz	�������9�e������T��ؗ#��y�z��`��c�Y3p�V��P~��gVj���R21|���j�K���-��|?�{!������FB�hn�$M[Ns�m�t� 5��3��t�����l�a�<��t_��O�S{��צ����@6�q�zh���ޛ�q:���gԽ�{�y�lУ�-N���{�m�^Ύv��:��o�����f�6q�Q�����M(�)0ӈ䉹�х�D����-���`��l]��N|�?G�;��3�V�i@a����UY{�A�F���c�C s���nM␆���(!�e�gx~�ş��y����-�D�ޕfY\v�@�3)�n��B��CPBT��)fh4!��]�t�A�E�Iq+�?
C������m�>xTl:X��8v�'��E�"�3�I4u2F+	�A+�s��r3�䚴������Y΃�1�]&����v���j���:H_a��禜z#�$�q{Z�P.fY���������C�-s^d��p�A��9�=����<>�ݷ�Bm��%��Q;z���1Ҟ�7��~��P�υ�xG�I����Ca���g�w��J�Ԣ�FE/��)P�Q��JJ�����@���_/ܣi���ܸa�6���%�0 Y��H����^K����/�[1Zs�@��v�Y���JX�G�$/tF�y��+��D����?� 3T+S�Gs<x��_�L��l��&k�5�5 ��?�-�t~]��b�~������&Pc�'��0�Y�Il����u��䄲)ITV��y�R�/���r5�@U�v��Y���ю�P���m۬�(�������BtC,V�Ssa����<YO�k2Ef�Sg-���+��=�Z�M�6
�j|d`��{���ZoK%,[�4J�L�k��x��Lw'��_+u�(�^Wҏ �JWm�Fܜ�%� �gbRFV���/,s��Mx�~�g���A�&U��G�BV����Ƌ�PDMQ��mn��߬�n. 
�&����!���~�C�pԞ܉�*�1I�I�.����ܼIltW�H*>	���k���@W�����R���V_�.���@J'4p>(Ɓ��7o-�񛡶� ��4Q�>(ޙ�V1�YK/��~m}�H�2�[^(��IY(7���~
�������}
�O�NJ�r���u�\˶�Њ��M�Q~���oUW�`��}c�j�V�	q��En�֫jFhBl򅶍4�;[n��;N����5՜f�C��U�
V��OI���-��"b���6��Tlfցd/�vFr0��\[:����9���4Z���Dn��_��!�ڮ˶��l�d�#�$�"�o����M.��&�f�����Pj�8�4�HS�Cr�	�p�A�kǲR�l��� �2Њ/C8ݡ�9A;������#O\i���nF�R�Nۿ)_��T���➟.� 75)��*Z?��a�B�����@iA��_5�5at1��b��)� t=U�X����XCW3I��I�!�.���U�BGJ*�d�2/�u,�m�,i���|�x�9ߙ}T�}�հ����dݱ!��#v+h\�60R0Z��ȅ��@���7]�,C�W����L�L�1b�p���R1It&Y�����_2�p`3\��D
�D��E���&�ׅ_U���Ê���eZ�M�@�l���(g�������/h����1ϟ� �s���0-8���5w���-����S�v&���T��6�|�34�V�)���Q�ϡ��-3�r�����a��-h~~e�g`�iHc-MKRߔ����PS��<�_BS�8��]FA��N�]���T�E3dO.��ģåꌞXώ���u�t�7�{� ��2����_�k���qH���%`����s{�X�� < �����A������^"�\D��� �'�p�W�p�u��q"8�((\ÜMގ�d#���,��
E51�2l���ڣ�wt£I�+�0��*A���
�� ��-i~�~�q��4Ǣ�݋)�|p�2%�FH-Rs	��k�X_��K��e��@�Q���ce}��ޯ.�zŨSdR[���=��<ֺfi�D���y�FT1`�5]���x��Q~+X��#������i� ��M��MhA��M%�Y�i�+�����W���s��;�/cᣊEVb,�KoJw/���{O�i�>Z��� 5����z�g[w�e���jN��1�l�a8�]E��jt3=�t�	j�������W�������ğ[� ��L�0�_�t�����=����n�rt�%l����v=qg�)�� �j{�9�C�:̵�����#���z������<c�jª!�r����#k6 Ph�������>�C��*v��p�`B�� bA��\ݡ�t�ҍx����5���J�}��$X���G:���D�*����6�'�3�`97����[�"4��.��y���HObB4_����	s>:����G��M��q9Vn����[[ۈtY���T�z�G�T}"�i�0�Z�"t,�[�����@��-����[��<���"u対� �J��m��h%`%�I����
nΈ��̈D�Ț�������嬁���)���z�vI���Vb�X�/l�wEL�(Fo�:�N��΢�42-#�:�[�:S �N]'���oLISֿ��*�)����wH(Q�nF ���d.���`�qڟKX{��(PJ.�hM���6a\92�/a�F����xܠ��Y<��ϐN�Қ�˘򰦾o�����N9��-.@�e��HBH���9<g�O�[�����t��ى�'-aϜ{���؁��X�����d���>�F���`i�P�m��MR��3n@�p���4d��G�s��4��C;���LAD̔�a����rb���Wz� �nUbG#�/{�&������z=^��֍��05$mw`Z���w��N<.1I��*���a:R�ɽ՘��p��C�X1$�����3C��,��@��|,a2΀z�`PK�?�OZ�'���r���I`ͱ�ѨX٫|�i�%�r�l�&�ivF�cֆ����ك��E��IyH��?��#ٙX��La���~g� �<Y�ș�<dS)6�~�@ϖ�35O_�,�⠍y�Ѩ!�0�0��T�2Ϡ��,�H��r�GV�+��M\�W���cg�˟@�������b�	�g�dW�gr�V�rwB�"��-�����v�s0�^�0��+|�bԵW���;���c�+n�m��d�ZKW�v�����)V��aO��]*#h��]h{�m0�>%�%0���jf�6+N"��m����N�"��V�4������wD��!z�@g��h��-6�/n��n�ț� ��J��򶙴
�#�r�LXs?��J�3���\W?��u5ߪ��wࡧ�s�s6�S�g
������д{�nK�N��W- �r���Ee�,*��(Ɨf	���F��nt4>��m���^�U�4GV�zu��x
X���x4�qί�rF�Dd[H���K�z��OXm�f��B�¬
+�]�.rGHդ��62kɑE�c"EdTV,��O���%�I������D�c�Q�
�=�C)up�
�xg�Ϫ"���{��A���8$Y�	�~�m1�
������{��AblJlL�Ooc�n�8�����#ϡ�U��)�q{	d�0_?�5AkD�۷tC��V�������sH��V�l��&�"l�b�*�Q4�j���[���j�e��V�Y���ټ�b׽�`�!˼DO���Z��H����W~^����Q�u1X
�����q���v=�2���A��Y�-$9�+ő�l�T�h�&��]*�>.Pv�N8z_��=j褻���5�]w�/���t-�-�:;,�+����^]~	�++p�;�
�w����l���E����_�i�I�"�Uk|���~۠sI�DM�e�뵄"+��*�_i,P�!���aO��|"0ޓL�d��#]����ܼ���y���n�����8q�%N6��e�~�Z'A���N�'���H�/�`8���ɯe_/i�G'��_�&��e�y����A���Yшr/5��|�1�0��5�:i��+-ueL�yÖ7�^e��v���*��4P�w�mf�у���3��;�sz�ѻ���7��
\@+E�ˀS��������G��d��oKe�Z���T���_tkKx�ШP\�e���52%'Q(:�"�����O��<^�2�F�x!h�s
���c���EL�#�KP}�:�<#��!�)+�(qݐ�2�}/�1�����*&-j)H�"��>�F��q�M�Q����s^�p�@��@:������8u�a/�W/�>-��o
Q2C��L�}j��2\fC������~���(�Z�^Ɵ��^e��m�L��e%iIK�����!vրrw=t�҅��'|��
�o�!�y"������ ] mz�����k㗛�����{�7���O�Xш�����԰[�H��9H��s��s��?��Q\̻m��-k@Yu��Z�����9�� ��3[����iEx�cΕ$�o?��gN��n~�b](���Thо�m�ք�+�x7�a�4i���Q:�� ��%��#��k���|ad%#�����$X*�4�v0v��a�A�ڕ�xr^9�~��dp�u=����S�.|�飛�h�鑼����[L�5E��	���"�ɨ��{���c�~#D/��,A�7lh���E
ti.q7䁽�+y��'��!�ZH���~5�e/�9�J�B���NH
�呔9�g _�ݘsNu���s��@�~WB)��
kU3xϞ��[8�%|�~1�n��/p�t�m�#��V%Q�83�̿c:Ԏ� �e�����m�s �G?� J/�3�m,	��m���d'��N=�[�P�	���Z�i�(�dӹ�tԒ����wIl�2���g��9�@�$��分�S��'W���_s���DQ�����4���	��՟��O.�"{��~�C4<����K��P:%J�;�%�̓��Ȍ�=]�
�w��f�5���&}����e��\|T�}�����K�*����w. �H (��н�����f�V]=JQ�O74 �p_��繅�G���Y�H iv�h�S��!&r���q�����o��	��)�_w6V5l�����BW���$N=�%��~?�`oU'V����K�D�v��%K=iN��\�C�0��Ъ��O�jeiq:�Xl9z�L���T�,;��t(>[��Ԛ:�;i���M���J��S;�a݆�e�[h6£�IX� !�x�#����C�i+��g��l�Q#%�g�� �X�"B_#��hи���n�us�|����M�DA�ҵ6l��r��a�v����>���Q��n*
j)8K�O[HȮ���<�h�Z`,_�$������!��o	�Hܥ�x��ڝJ�#W�S\_����A^�����z� z����Ґ������#RV�x�P�X�<�� �G�h�6v��ȑ�����B�G�]��ˬ��Fx���]�K+54(I-�teRlX�ԎB�K�!��\z5P�݃�5x��Ђ��<=��a��bE����զ�zG�?w��Y+�SQ�����S�-�ĺ�rϞ����${Vr��O��q�i����r���T��Բ��|3�%��^a��@O������y �l���։I�/ܞN?F-q��	�,�����	z�6����9W��*�̋��2��l������AuTb�Ew�\:���?��Y(+MFp��َ���B��l�N��cn��}���b�П6�j�>��H����iI����Eu����>Z���k�F;��%�Z�N�ᛘ̮������a�P?~�hE�A�Y�w?˼7��z��8HS�-� �p?�2��#V:�4����WJ[�1x��T�w��M�m���k����ԣ��}��^�ݫ��mN�eB����EAf��ӽ��&K�r�|�q��,b��\��c��3W}k�Fba]����%�E��$���l�K5ZE
��|������oUn�~��7�e^�k��N�{��D�+YL���֝Ǔ݉��C5Bj7�%g'-AsF�K�Ay��ن>0]���׽��^�O)����G*kd�y�Iy���-ws%|�iT�ƥaD ��7�$`�,�B��=Y�٤���r�\,dt�)�5�n�x�㜞�&�#���y
�mdLAXK5gt���Ŧ�Ya���)􆦸z�����U�}���1��Xy`k�2"��%;�M7��׌ZR���e;u0�CV,F���}���� �-��1)���E�'g6�_��*m�V~��5�;H��ϳkl~�Y�7��δ�ؘ5r�1)h��4ӝU�z��"�M}孢��r�l�>�/	SHʞ2"C�6�YX��5�&{�-Re~[!|/Yu]7\·����)V�FK:{ �o�~]�.G`wZ��6��\l�["ڑ�W�<�2)U�ұ�d	ϯԛv�XT��Y
��j<)��R����%��gS����a��)�L+7�ʑZo��B��e+$�Z��$0C�w�b�2us���j���Y�؊�w�YM���ž����L�B�/%�1fW+G�y�Ҕ'�����S�)܇Õ�[\�̒���R#X���y�R"Q|I�(�Z?� ����y	[އʍ�AcP�.'j5�3�w.�ּ�.���bvQ�ݰ!�m�3<�&Y;���#~�P�.�J��b�u�~���2�,O\Nhq��]�4�xY���㭛�A�%�9wUSl֎L�����s����U��EI����>e�`��p|w-aS�D�uL!Kݤl/�{��U���B���4F߭lg1Ƶ�m�"��]��O� JH��[�Z���:<�W���96��h�K�Z�x�@�k
}�G��or{a�H3Ԫ��AK˟M;B8s��p���(��5�(9���,*tco]
M�{�:���-~kg~�C
��A
�
j�ͪ����(%99��F�"�3���I@U?x6��\�j�c�&pi`h�CG^�����B$F��SK"��[f/��ù;��r��`}N�#�9�a�RT�<x�
5�
r;��^a������"�)�MO�ٵ�����o!(t'�1M���J@�� 5n�	M��N�����v�2M�ҜGz��2��ek?c�12v��V/th���<Lm�'v3�G+��"�:�a��WR$�W}d���Z����=FP�op�1(֡�yp̀9�Z�0�-G�v�|5��o=�R�0)O�1�F�+�R\u�oz� �5 �^�'���ˈ�o!ˠ$l@�\�ܽ�������e@��~e��� ��'��~�k?��?:��v����e�J�z�#��Ҹ�_JJ\��$F���3~���HU֋��[�a m�g��%Cu��K��t;���`�Θ�T�������� lΦ SJV�vrcc��^O�J0)�Q��i�m �&4:�]��y��	%�� �:1V�����'�W��	��.��yBTѽ�.��+���6>EyUɀ/J��w�
��r�������#���<��`�lA8�x#�X:,�)����}z���U��n���G!0��f�Bv��n��e��Z�g��
��\��,�gS�R�>h�5 Yƙ2�A�I�`�+#�v��gd��MrP@~��÷ݵ�j����K���5r�U��Jt'�.&�X�p��;�w<���Gj���+,TZc�{��s���x�ԑ&zY�V��ar<�!6�UI!����T7�{u�3��j`1�����2�}!d~z���W���eĐ�u�_��Q��}�k��r��߯��A�W܏E4|X
o&[�!���}G��%��	��mԆ��sKټ�,��w��$��._o�P�hGy��K;f9��'�A�����3Ca%R���<���e��)����)7�l#�j�s�bc�E��ʩ�^�b��v�>�ݙ�w���A�5u��L�[�����������f��|GUo�\�X+%<,��$,N��kC�}F��ŗ��^���>�����t������tƆK榺���g]��E���̀��q�X7+�����h��+���ҙ\Nn�Y+Y�(�U�(r��/ q�����e^�_D���i��mY4=�����2��`2g�x�֒Q>��bG������8�OŁX�$^�r�֗˩]
7�;�R~$ۮ1�>Q�o�띜�~F���n�,��B���#�D�[msǀ�^��6���mS>{F���M���(:J��
�d�_
��͕i�s�/�A���Ȝ�����ܳs�| t��I�����0��Ͱ�{��,��C/{D����U�A�Y�G����B� 袒v���r�?�8��
�
�\ �p�b�T��;��Z9\�
XזL&6	o_�:'-с�yI���m��	� z�P����wE�M�m��0���u�
��V�� @&�PUd��渕�d�JJj�z�o�||���]/C�h�}+g���Ɠ,6���,���RH.����ԅ�.ifL����,[r���CH�hJ������y;�ک`D�r����/�պ:�����E���DQ)���<��R{�k����^���l#n��"�T��zL�rܚ���S�K�ʭLɶ>�Nc^��t��n�ZT���/��#�$m�X��v�@D��%]|���EEФ��Q�x�F����a5����{�t"��Ν��6���&cG�
_�#���A����F��LB}�k�(����E���,GOW-����K�X���̕h�s{��⤟<LXը(�N>�!M2��Y��qq�A�j|h(`V"(�bM�3�I�#��_�S�a�	/�-E	���1���
:�kW<4��<����U�<ɑpn���Yή�:1�&��:�����ܦ�;����N�g�%CJ�߿�:� �_�����~���,>�(^jҦ�g�'��?�@���B���Q�U��$��sK��@�,�m���m�|.��S)wԞ��C�6��i����bը�$� ]QD(��N�O���o@UA��'��Ӗ��қ���(��*h�¾��ĊPѼmm��K��O�'���-�����l�o�j�wH�I�o�	c��m@
�R��o���xQ��o�����[{��>���4<�&�m��3���XcZ�.������"U�gqa�)�k��Eh�Jv!�b�С�p�[���1��'�C�f�@�+Z�eR�j$��g�g�^
��o/=澵,�b��Īӏ�e��C�w2L�|ǧI����m6��it����w�oM�����+t�jL(.%�|8���\�)ωBd��;汈�8q1	� ���.#�)�w���t� ���bd����� ���	�'���8�5���։�P����ˡ�	�a�E'�ċ|�`��M�Iŏ"s�@<h��d�:�6ƪ)�FU�/`���[�@�>�gČ���w��܅<$��t��9/�y�b%:v�3�K�6�g�xc	�h*e���A~KV�`ζ��F~S��%�p���I��'-��:�n(tM�j�ڔ�w[)�j&�h���w��3C��at�d�]�)��J&,�t��q���Υ�4�wG�)�؊�[�t��_ �?��FU��锴����<���1���40gU�
A�w��-��p|4H 3B�\4�(��ª�Y�Qї�@�T&���(`\y��ZOȭE�k.h-�zR!{^�\7g�XJ�N<��^f�e����J�����,�P�M�%�Q����T��M���΅e~��s����^���?��aE�GɌ�w�2EWŜ$���Z�e�~�6-r,��$�Tă��U%�E |��L�V7�1�L�߉ ٴ��"��G_&�¤͔}�Y����ma]�IY�U����,���!V1$��8��C<af�+M}��V��yU����p�A���	��:����t	Y_��1��ȃ�����Lg�� ;w|�c�h`�s a_쯡�In�A���zp4�YC�2�y�J�u�5-]��8�=�U)h�~���m��-�4a�N7��o؈&����0m����~,g������
@0��r $+��[��be>�b�� Y]��H�֢�ح^z-m3"��w>��R0��	�FH!��.a~�8��2�}@�Z����a�,�zN�+��|�M
��J�H؋�,��3N��*ˡ7�|��k�AG��R{��V����"+���~���7��Yì��*��Y��wsm+J��'N�D1�aπ+m�P+�4nϜm&��mM%?m��Y��ɽL@(�:��8��-�	��Ck����{^N
i����:2�SǗ�P_įO)�WW�1Ph��w	���/��v�������(K���z|���J��c�0� \���r)AW4С:2������T�,�Nhf;g�VAv�����(�H�z3���Y�8sP�w�.V@Ơ9���CĀ�d%/e#�Q�(��J����x�,�q�a3�e�-��$v`|é�F����<� ��~+N$� �����cV��p*L�JT9'0վ�V���������	�
�|Q��ґ�����	�މw����#���2i���o;�^E�����%��x�s���U��yA��x�"{���'�Jy(�������b3t���e�.�����|� ���>�QV�A�O�,�I=�;���a#Ȣ:Ծ������a"�����j��k����a����8��O��ͽ}��L@�����R���q�'�Z`�[S<;=�'mh�M�����Ab�t��)j��a'��[웫�c*Y �g?����c�[
��H���%�Z&��/�C���Ⱦ��^�~��m4�G!������2<�I$�k-<ݝ�ڿ!��KLPPí
b��|��Mx=ܽw]9I3�H@:������%v��*m~���d�T��vMY�S4}�ER���@]i6h��@�L��
����;:]A���˱���U����
��-���z7~��v�0W:KYM��r�Q���ڛ�Z%Hd��>{�����V<w��A�<�Wfu٧2�"��������?⃉��Ά,N����=]��R���u
BO��%�J"� �K�_�N�N���q���`�;����K��
TQ�__^'��S�(k3vJ��[��4KH����K(�2.Rsf4������n�FM�R)�Q"H��d~��K��z�K��|�f���`+
I���Ȥ�Re�����,"B򨟴钤lر0<�&Ot���ѐBc�%e�[fI�um�l�(]ݴ�!�j���*I����IRw�xb׭����x;��svϥ"O�,�V�4 V��(ҟ�X[��6�i�]y����z�B���4�6�u�׏q;�w%�NC��)SzH?c��w�!��=d��N~�*'W��Dm�MO��.��3f�H�A�W��o@h��ْx@|>I.�l�n��|�
�����~������M6F4}#�5՜�܅$	�$���p�qc)4�p�%����Z{)3�	�~`}B+���9�c5$�e�w ٛ�G�NV�W�ŏl)�f���m7���#L<��7�|$hX�M�D�k�_�����ZB�_���-��<ȄA''���YG�b�YI2�4��R1\�gB��8���tU�����Ҟy�:���ɛ�Y1�F��\A�]��Z��tֺ?
u����7¿"C�C�kJ��jK��+`X�Ӓ�(6���H	���͈Ⱥ��O�>���F���4 ��[���u�*^v�����O�V2�6�e�Ń	�D����S����紗���)�Z���|�4����š���`��i�M`�G�CL��p��iP������:2����V���D�y�-�ޱ���XƐ^�n�-A);�Dx�^�:�C�X�@�1��?9R�Z_�Њ���J�D<n�_6ٍ!X4����&�o_f�)de�]���P�~x�|�:,�� 쳔�&��r^���t�Ia��� �ڏ��� ���z�]�8��|!X�#N��;�RH�e�
��^�0�j�[���b�d
�0Z2F�G���Z����F��{��*x6^[B�ۤn��al��곦�����i�y�q�7��=�����i��B���@ �("�5ęqb�jvej'�)^�
�sD�7��I,0gzwy��;���¶^g粨La��7�:��o������\��Y88��j����S��F�Y�ժ��6����i�? BE�b���l�.�}���Q6XI̗Fw�P��L��C��o���-�O�r�<�9
�3<zW9��ۼ��d��d�ko}��LM|	:��s'Ս�����[FiL�%vE�ޠ�h[½�Ϯ��p�!�Vb�Lar��'ّ5_��V�P�Qަ��Ze	��q[ʴ�H���,24�s�f��&1��_su.(���&�),̄�g+@%.8A�A�����d�.�i�� ,dPdow*9x�oq7�;]�,�NX�)dĎ��/O>�E�tVdwT�Dj���֖��I����^�"���(@̧�~��y��Vx�+MW;�6 �޶�Aw(�S�Y�q�� `M�'mPxW���91��~/x͝���i��w?�?O�>'f$�6+txU��\�N���$V�o�]�ɜ�h�F��۟���_
�\��J>Xr d�4�����6��r8v�gԘ�V�����T��ֲ'�����{�&��Oy��5X$Y�IZ��y�y\��Q��M3�����s��P9��1cask(���c�.�\�J�	�l�â`��>�8���X9;�=�X�D�CU��ŖxZ����m�>�z�z&����Ώ&4TRbRYU��obi5���Q��[N�)֧�~@�j������1�n�{h�L3��:$	�VH�]b�Ōu�.�5���>��g����|tl ������Y(�X�S�UZ�w��y�K����Cn���l�o�\��m��%x1�i�"MM���*���:���ʾ%�t4�Z[��+�Ɲ�/�㞸��R7�bF7Ӡ�?����1�72��^�"ۣ����dS���гNL�ʖ�S��q7�@3w��
����-�_�Vdr{x�z�\u�s�����u���}��^x�ʈ��(�BVq��mۓ�~
���[�E�q3k�xr�dי�*p���j盎Jq	X�K�R�B�b�,+)���3���Atmm#��I��"��w�-�!��;Z�!h��'��v9��8�	�0il'�9+����H�hKt9��;C8T�җ�������CJ����7R��]4ƟaB��jf:��Ť/lH�����E��W�T�^����/Cl�xg���|01�U��c���#}�+�
��L7��{��+s����7�3�Y�U��7,d�Q�^8�*�q ���XcV<=�L��n�ì�PyR����P�[{$I�i�#�z!�ń��2���qHTNÛ�J�� Ch���e�B���nF��UnQ����<a��󠘳�c���g��0�М3�K_*��y��<�_0c�$�<!���K0�@d�	%��0���q�Љu|V�+�#�f�;\�E]����٫ hضʜ~�������g���XзH�=�7�en���<}Ʀ�t���A���9VA�Ke�o�!Ps�TT�\TO'�m����N� Xǝ�m��s/1����ma��Ο�6(ĩ�w���t�O����?7�D�#�!8����ZOƺ��g����ΐ��G=���A=�.(�{G�t��h-{_�A�Ա�����*u%٤p������`�m��Q�Ea���8�q�A!>Ή���b'י4;H*9���u׭R��L��ksqRI1�_�E,d7=8�
���K����QP82�r2:�b5�b��A�M����=�ԧ��B��s��}�=�Ս`��j���z���y/�W��u��+�x����@wh��^x��8�"7->ʛ������zeO<x��Z"�+_�����,<���3}M���c��i՚����}d)p��c���dA���</�!<�8:B�GV&����=�vJ�lZ���ÔEP�Ξ�?(h�9t���\#gj#r�~꤄`�-�2��g��n�P
dޯ&��垆%Î��l}ܱL��'�Oi��ڤ;K��:'����W�C\�]�.;4v��|H���S���E>kIz�*d�R��v6O���$�e4/�����(瘴s a�7)A�z�!�����Φ�D�s<��U�" л�X�8`OG=Xʷ0�8��=5	�}����wf��Wh�Ǝ�Oսm �������a�gjp����f~�}_<���<�u�����6�|��qL~���{�ý}���S�D�3F���,��#��|�c��U�S�;IP�+���$q�1Um��׳j��+C�ƕ�&��È��PK�%i�K�6�C�l�� *[5�h�,xCe<�Zn��&�(F؆���(A�75/���EhvE�-�
�7�J/�ߖ� 
���oR��Q�&���YL�:.,W�S$�3!M�|*m�����0���D/�˰?�)��Jos#�K��>��Ʌ�>�;ʞ3��%U�~�ש�JN�2�Z�Oe��=�hx��XfN�}�/q���?��8��"���P�骿���͠�u�6���A�\�ȴ	KL#���1�,��Q�@Q�E�>#!V^��L�s��2ɚ��ʮ�_��8�u&����Η~�9�����嚧V�fc�e��lD��\]H�sע��
z�❋�����:�?�5�uZ��Nvl�9��S�S���l;���q�b���z�Τ[<Խ��)�cH�����t>F���^SX}�%Z)��}*M�[9k�ϧ���m���#QO��~6΍�O��g��J�ύ.�q�������$�3�hi0�7�^��X�R�(���\`(xE�e����U�kd��.le�<i��ޕ�<�$�
��?�!r�b킶�
���s�/f� ��|K���������y�����o}q�ɲ�p�G>� !����@��He~�<�9�~���(��X3<U�m�'�Xy���x��_��8������/n܈PQR�i|���m�7_�^�y��x�O4�Ȯ��wMg��b�����v�5OB�˰��{qD>��;l%�ܝ����d���F�z�$��چm�2ܖ�[{v���T� TOZf�)��'�?�{(��,T������}PFcR�:9���Śs��|\�O%�����%��&[�?�Zi4T�����1�^�S�$��M�(��r��$�����L���{h�5�D�|8�%R�y���)�Ym
���Y�	�4�A�N]��N>�Bvz1�i�D�@=;p�YЃ"�����MW�i���HI?�w�2����RYz��*��z�\����F[�)j�hֺ�@r��@G�5�����es��r&Pa�Hl�G�K2U3�'��9��:v�f����S%X���|��b�7������'�'��'�lʡ/���}H���J�[Ls�2��
���;
ZZ��y+2Rֆ���O���g�4I(�U�K??Ɉ�$����+D�9���#�V?	I|	y�����2U�-�㴵&�f��|%-u.��3ζ���&2 �?+w���c(�Z?��0���d�7�|��ޕ��=/�YHZ��x�']=�|��&�jH�ݤd<.d��F:�'vRk}4��`�����8�~������K�q|h�`��N�_qP��н������Jn0ͩ�)�s�Ce2(�ˠ2��0���� Ո�c�W$��r���~���U�^éIӟ�Vk�<@�D�w|_�ĝ��|�f��Ŀ[#t�󞾓_<�B)�MS�b%�R��p�S%ЅD��H�$r���d��e7ߟwkp�twV��Q{-�{
��Pq;4L��j���\�(�/_u�PU��P󪑦?΁1�ԪwS�g3�^��Ib�"ϳ{f�AП��$������g8Ks�,�ǭC��/��k[`���7��)Z��r�fjx���>0v�ߵs__�~ u�Be1�L5�M��n�^���hN�ǳ��t���`^n�X��p�-����k�{��i+怄Z����Q}s��p���(g���O���V[��	L��汧���|j��H'�����a~���!�U���'fSA���m������,�_Pf�x4?��ʴkSkڒ�-a��f����ΡN2M\�P1��դ�Z�W�5��l��$g�f(�͜�u�������<v����&^u.�ha��x���k�����#�����m��m�Ѭ� eu�c_�P�L�����_>z|�"鰄�i�;�gU��9L�Z��Z�<��/ڎ���ƲUf�>��SR��ߟO��>h%��-H�����H��g`s��� ��}c`Kg��?��M��t�����,���U+�2=���y����Yf�U���B|�.�U������j� �@.P'($����ϥO:s~J�E�\�\oU�=C�>!ʱ�>˄�4}+�N/\��gt��!�UY}D�b�f�3v�n=��x1�<2�[��lc��9�6`�5�8�[PN�:��?&"1���ذ������˯)#�m���m��6���k� oK�)_a���5YhM���h4r.�J�/�I$��oЧ�P/j�?봪r�Z7�!4[2n̘:�4��\��!��WG0ƌ63�~��F���6��JQgsX�U/ܪwd�`E7��ƻ�
���}���R2�)v+�����g��]���b��Y����L�1��f�,�?I@g�(r�c��3�s���J�C��T<ե:8Ν%�V[�������6f����,�q�>d� ��[���lj����WC���)ަ	ESkO!k�UJb�=L}Dqn,�f}c����grZ��e��A�;b�5<;�H��Zj�E\��?�:�w�}�tV5M�-�/��&sf��G�K�ך͋�N�sj���T�E^sh�E�3 l�U�@k�>��$�jG+0}���X��0�fG���=S�����H�)N6X����7~{b��7k׀��y9���q*C��~������F��J��Y�Ȗ�Y �Y-�s�LC8���t_��4r�Z3'^���^������K^ #g�բl��u�Hw3�U%�>�l�j&�1lԩ��j|�p��6�ѷǺ�)���͔��;(9HՋ[!���kz��T�+0�Z�.���1�Z�+��	�JJ-Q�]���c^��t		��BSc�lheM�0^ 1^��բ���K�;ې#���ۮ/�
�Z:n�	�7�-������2v���X�o�q�~�E�C����V�'P˄��۱�\�SN���Ke���}Aξ������Kr�N��I��@�N@c����4�)�����	��C�q����ݛ����{���]TY��\0��]<�ꦪ���!`~��E�M�l��P*�+��`�%��ls�5�)�Sh��]1��vo���Jz�m�3
'��F,�;D����kU��p�ز���Сt+���ɀ4U��>����&(Y���U�Ӧ {|���17OLۄK�R�u]Z�A:�Ȗ(H�Zp!�Eʊ�蜋8���O'�m�+W����>|PN߅cҀN
]�����i�P�Q`�����̔��EdM]0�/�.�r�Ǆ�,,me����p	2�����r��N,�Vz<���vO~%��c[��]�a�a��������j��2
��,B�Z@�'~�,}��u~TБO�#�S�I�x�X�j����d�e}\���3 U�������q�@���1�NU����������ƋIrٓ���%\�
쳁��xS7�N3l�89�SC���M˳������M�\��P/�w���.~Z"�5K���lD Rܖ����r�3��bZ&:x_01L#MA�x,�-<	�o�I�Ê�o'l��f�g�z�u����od}^�Ĵ�w�/����b2�_�yes���z$��=u_V�ĝ���*|�uf����W)f�U`ҏ2~�u�z�
4�˸��K��i���X7��h��EK$���v�E�I7��ð~�H}sy��0ڃ���:�����
�}Z�n�(�X|���wWv��w|J@����~���g/z�j)���9Jܧ�Ş�ˢ���vשfo���ˬ?l#oai3ŀI��n��xRn����̂Ƚ"H㤪�,4s%��|���ݿY�;m#���@������ivj#�z��Fdm�Ɓ2�����	u�>�	9�Ձ�
d�T�
�Z�5u�_���jΫ�ԅ5R ����l}�4�E<��kG�d0tr�D�PS��E�������Ԉ�Q��xYw�[�6��n( ��^i���ų���q��4�W��4��x,�027��N�`u�pK��z8,�8s���vn�~t���j-G�]�5X�����{��`%�-�>g#��e{���@�S������s���%�F;t?��}ᘈ�l�4k�s��x��dyR�7��ķΑh��Eu�,�'*�E�KGV�؛+[%N���e����L�����EV�7>��g�K�+�v�t�����T����Dz��6욗��ig��s_�!�^}`�2�ʘ�9�˘�*�����TRyt{�I�%��)�Hߢ �h���E�OZ�̣b���-6,;o �ٻ#�ZP|��bj�6���8���׍v�Q��ǅ΄���)!���᣼�ĸv��pg� .��TpՀ��ʳCW:s��$��Ơ��O�T�l�x��w�E��%<?[gj��̀��o8�L�!B�.�$1��suj��[q�"d�
̦e8V�k���B��T�(=B����h����/թ��Ƨ^���������0?��_. ��̿A�G�,�#n9�
1�x8�X��W�ߙ���**T¾��:�^mW�RJtپt��*շؚ>y�N�����	cn�����?���썳_ZM���)��$\��QA^4���xI�>?�][6Ռ`<Pԅ^|���8�X�9./.����j�\�ZP3�Cd 18���\�\rQ�R��u�پ�ރ�O�^[hM�x���w M����I�ь�A_& �(%�bS٫�tH�`q����j%��:�
Sؽ�S��r2��ƕ+���Z�/���@H:�N5��Q��E�=�E5��*��r���;�seNxD��cq$�4c'=�fq��>sq$A���*pT^��@oͩ�f-h86i���,����
���JC�u&2��m�4}��`�CS�f�2:���;;�rəĬ��������:hd\viemV$f�>����V?�:9>�O���I����e�>s������҄�(��Y'"%��7uS�$��Qļ�D��v�l������R���������;�y95I��4.h~��n�=5[L),嘾�9v��N?n���~&]]�!v�^1[��x}�5��'��S%T�+o��X�B���c� �} @�_9؇��֟`����)�T,��ϓ�}����-�F�ޏ3`Px�ct����
1��)��ϙ�U��r�z��ͨ��qQ�\�L/���
���бG��! �K���C��S��Q��-��a�G��E��� ��M��nۮë.<��]��s���t�����&���*��v��'���3sfŢ�Ox�ؿ�
�aO����V�*�-��R�>�� �(U�F�"N���`�Q�W��)�eZ��4�K7��7�(F+}�t��n��ݽ��M3P� ^x���m�]��ӱ����l�*���)��F����&C�c�(�S%f��20���iz�"�>��:2�{��լz�8<u�m�E,m0���"j����f.�=�`U�/�m8@��5��D�.Nr��N��UB����QC��rX	+�o��B�6�$��ۥ��C�S��h�03�!�S�_�9Brq���j�h�<VY��$T��Ew�н��O��_���K@��Ǒ���F,�B�P���<���0��B�̆�k4�l��	���|��ɚ.rv���tmƏ�l�Ƞ	���&ʹ�&=E���'05�I
r�na�� �������$���Rgv�Ԫ/aD�O�}��u'���3և�6=�k��������H ��wcm@�,��Kj>�7��\�xL�� �Ţ�ާ.�&�������fh��ҹ4�jG�A%�f4t}������(V'H���́���`.�Vӹf^k��O�G'��ѩB��/"x���u������['�������U�I�y��/y�X�ʈ���i������K^�r����)��������|�2�|�j!:uzj��6����F�;��`�h6�`KY���(,�B�w�~Յ7@)�U���9*%.�G�� �b"�"��Y.���򗰱��$��KP�q�q��.��IO��Q��Z�}���z���Ġ�3u�[�����mc�c�v|�ʮ��=��舶7�ܼe�n�9N���)�%�#�,�q�a�_ks���>�U�x�s{%bS���X7�G�rƊY�+� CG��WK��U��i�����;�^9ב{QbG2�7�i�_�A<+��N�襋�H
2	���4r~�SM�ߙ�+��e����b3-���&\[��ϙj�S���k`��VN��1CL�J�C�
�N�PI�Mα�V&�iC�sM�Y�F������������B��ez�>�ʲ��!�� �kv�Paw �֣�b�oK��aj\B�h���#p�.w�T�إ�'r���n�J P����2a�{W�\��Z�lO���h$�0q>���JT��S�{�J(�"H����w�7c!���x�>L�Z�'"2^ob��,�7�8��,���qV�Rيnk���-�<�^��p(�#X��%��� �wQ(&-�&������=E�&����(�)���*
�x3Kj|�j�
ޠ]����-\�R�5:Ǔ�m�W Ք�� �J�7�������&agf�+���%����Jڛs�j�!4+���e�h˕��"zu1d�3<FJb"�9��X�A��ZB@�۾+��s�9_Eߏ� ץ�a.���WIǛ�HHb���u$A��ż��}��]�yf��o�������?�Y�3�I�]��ős��׏툋���C��lnl�X���T=0����s��"�|���Q�^c/���y���]���D��s~*�H�qG���?�[8}b7�	F5:u�
�۠H��@���ܙ,�nuQxzZ�V �m��qs��T>1�Z�����s@����M���\ wǫ��I+�� �&�m��	�D�����h Jh|S/�ÞV_v����忍;����ȧ3tر�;��q�>ͧ�6��km�#��hQj*�mW��Cz`S'Z�}:�m�,ߪu�.<�G8���+z�_�T�W��_^�LĪ�%���[���0i�E����ReR`%[���qf���; �&
3+b�Tf�Y:��n����^�ی��7i��0���f^7h�$o�g� c�eN����<x�f��p���qP�y�L1����	�q\������
�{�^�Rm��>6_�[h�9��'!��x�7���Z{�R��|dI��z� na�dG�}5��Q�~�?f�V�/6��⳦�]mK�$ �I����Ac��"����5X*`�#�ȧ�Gn��TtÓSo��nUN+��̅���B�~�i��ZLaf�*?y�,��kD���Ml����R("�H����iŽ���
�#�*T��{m���:����)�C�k���=�[�>�	�Of�Li��8Y��Hh������|�D|�\���Un2P���޷�S�W��碟"-���Z``���nX�oIi ;$ǩ�kE(��|	ϓ������BwD�+���\�j'H�nQ��BW�):���Y�[d���/���7)~'Z��q�J����ϐ䲭|4��L�!���ҽb?�a��׫���gZ�\q��˶�P�֖	����XdФw��Y��E�-Z{1��
(p���
���MCѯgޮL,��l�:�.�Qe^�/����B*����;���!��Q�*>��l������r7�,>^d��Z�+�ȱ{
��|_�4QjH��P�Ԧ�� ����<��P��*{�gה�{k@J̀�!�^��Gh� En�g TmcE�$���Njաn��{d�$i��2ih�4�5KCG�6ރC��BlE2������ݰl@S��<+�p /[؟��sgRg�,���?#\V�0����``�M�‗f����݀��.,�A�i��*�6���0i��,v�pr���͂��>�f*�\!��T�{��P'�����GI%*��I �W��`,&G <.쨏�3]�t:��R'L��Y��!5%�)�+���o'���QU\�CG߹���]ϡ ��"ٟ�|��_�.�?[��h"R]ޔ����`�}I%�{C��n�$�(�⤋}�~5�9�2�f�V�9k���ӳu�*�f�gQS�c��]�\5E��v���+�.WZ������K��nv�<��	?B�|q73.I������n|��/�s$z۩p���aT^����o��ö���s�<N��tjM�5_j(��0�������.��e�p6�;�c'���)�<X?����&qj���y{1Ө��YO�s򳙇*�������-��_�N��f��T�p�8�K!H� %��RQ,8�!�WxIːYMݼGp�RjdÈOCFx�%�_d��|x��2?{E��l@{O�������N^����j�0K��f.w���3���LD��A�V�������Sр@LAӬi`�GG5KE�o��}���q�1>8�ކ�-���pR�=�*�n�)��ֵq.�������#'T������ a1=��&"�kT3+��r�Ƚ���ϫ���9�\�6���[H�n@|u�/3��to�,���\w;~���h�3���nK��0;�s�[��C�$$���F��&�%M9⌉i�0a3�ՙ�7�ט!�b������ft6�6ʛ<���2��rY�/.����.��&�F�.zQ���`��̑�����V=��� Œ�OW:���S� ��M��N��4BFmh�����
�p`����Lb���V�ׁ5Al����4Sy�_f(��FΉty���E(��%wdg[�ܱ�َ���A�,�mӲx�y[;�ƾ�y�;�p� \NTa �N�i����а?0��0�nBOq�Bq��pzzҖ��QVr0ZGW��H4d��,O���p�3{L�r_䤶�\�"O!|�e�c��O�)�2�`��4�c�(i�ήmU�w�Y�ϾZwz[���ߴG>�8���5RC��l���z�Q=�
�E�v�;3w7�b���fH=�����]u����8U�ʌ�s����+}d��ଶ�Q:j���Ĳd��s+�x!�}ςj �w�� ����P��g��_Ζ4@�������-�8�{5��|SD������ň۰
v�K�NK���/D&�9�:�Y���ܘ��h���蟀k!����i��bKB�_a��F��X-y"���2X�(�K<�4�&F��%��ee�H�I�W�X}��i�u]�8^E 4ۘsm���L��p��n�9lW���rXn�?�ڙ�E"j2y�fʦ������ZF�5옐:	�� �D��Y�`Ww���c,�o.n��e���߶�4[�b��	\�[#��n�]l
ԗX�!\�$I�O���~Ǖ{Qkd����p�<K��������g� \j(�$*P7�?k
�������۝��A<�8W����*��ǔ�É�l�i���te;
��^�wR��3��zi��!��jlЫ�:��;j2��mM��fh��,�3!�Siq@��������KlAHg�I-���g�n� ��f��d�9"h�����N���)�6���cׂa�$����]FԵG�BC͹�F�͈���P�_���a�n���3b���������yWɊ�К�L9�H!���Cp{�	{�-��!d�A|.�Z>H�W$�%�4�z�.��5�x�?O���}vY�-�^��D`���/s7���kr���1cej��y)a2D�Z�4���G��}��L�"}w�������po�,	Wb�q<�?�ߵ���*�9�?����r�	�b)O��bhʌC�=x=�a�-����n���?:S�ߑV�|��2��(�o�b���?��ӞSʿw2���5=�HU��7��Г߻ԭx
,��5��}?ȑ��su���1x0���8$�ݒTZ�)��?�o%<����.A��,CJ }^�a�|>�3Ԝr� ����?�@k��������ؘ�,�*dнf>��3U��('���X���ܰ�Xj�E�Y׶n���@eì-����{�?����� ]�XCЦ��cV��k�`�U�_,�8k:l�CG�#8W,���D���e~`���K3�#�X�D�J�kOr�����U���%�a��I]����A�i\�>�Ρ��>5���(M q�Y
L�hdI��}�V�9�v��!�wB\� Z�tUQ%{��u.��L`��8�_�H��g�k��K�Y�N�S�h:���ޅ�>�Y1z�Z[m�\?2��QP���SZ�,cM
�P�L;M��E!_�����U���Іjgd]0w����e�� ?������e�la��_"Ҭ����%�2L�htH}I�ɟ��Љ���&�w-����_���fg$S3y�IqT	+��!��z��G������u�Ϊ���ܠ�)h�gM~|�N��� �тշx0�	�u�.A"SLa�����(��\�����f�c[�����7�vA˞�gj.�����E�T̍j�ߗ�}|O��<R�hg�c��zS��.Zq$YJ�ؿ�6�x�.��B�Y��<t ��@,���8�3��6��}����"�a�8!V
Z�����G��nf1k�bwX?2�srS�����v�پ�>��k_���c}=�U�Lx[܌/]eU��+��y�`��#�N�(��ݰ.h�f+��*#M9����������o��Sr��>�6�w���4�NWX�ǐ"��r@��;C�]Q�˜\�fJk��F���*HC���f����	��o9=[r1�M�a?Q8а��,��L�x��)*�
�=���:��Щ�+$B1H�M<y5����x_|9ꓙ$jE�w_�0(��%OF��P�c1�2�8�]��Z�Y�1H���=NwH�M��f�U�8 s���H_�N2����1����~p�[d5�A��N��4t�z��.�<i<�;�f.[�i\BDt���F���l]H*�&m�O���R���14QH����<ճ:>�m/��[á)���-�i��6�؜���E�τ�}��b�s��_�g�,�	R3:�R�HQb��Ԗ�_	��+�Ur��F�zǁ2�̼�Թ���M���}�txs|�*�n6l�y)2lY��!�ɍ�R߁�+�n�zW�!V6�Mk�o���t���hk�M��7!����"��T&�� &��ۆ-,$���_��r����]�$l��4�����A�k.G���B����O���&���>��q����t�v+���`y���,wc�z
.7��Dρ��;�z�����	�pT��H�E2ac����\R��#?���v��bf�ǥea&U����BaISoY�ʟ�zA�1�L&��� ��N��#���My�����!4�@�p]��^Tqw�4���Ԑ���Kٸ�/s�`"Dk�d㨁4Z5�R �r�� 2b$6FN_l�N�i�+�⮔oO�ɩO��t�����__=ǈ�`|��u���W��y��1��p�9f�AT�Z��8� ap��n+|Z	�UEG�Qj�s�#*Ƃ�w���~���왡��0��ڜ�3ش��[���z@�fң��Mk XA�jHi�+�S* Y PZ6�}`O|m��G�J��_�ؠ�����𥴯�ݓA��T�UV�K�+�	�$�k��{�a#��2d�Zp���+[�Q�o2c%��h���Z:�
.OvU�IXQ���8Ȅ���@~�5�jȱ��P���Rn-�k7��Ai0�U�[�Xuv�H>&�|z?�!v�Ml��%��R(Z�y ��<�T�LD0Mh?[��a��5��D�t��v��k�S��C�o,�{"��_���X4�ɼ�ej�_���o�C~���Ke��2!�v���#5r).ļ	,l:W������JƮ�76�}Yאݕ[��t��G÷���6}9���R�CHρ} LO�S72���`�r֎�I�1����d�ޗ�H�yʾ~���5��͆�#�[�XF�P��.U�Y?]��J�Az[��[�F@�؟y�Ƣ��?��w�b������i��f��_��0o�`�EG�F�"����oDGJ��Ӳ�J%�&���ӝ�$�G%�oW<@.�y `1W��?���`
Q>�<o���i�h�.&SH_D�R���������;�����~���ׄ���=��ڛA\y��0p�L�}��}�����0ec5�H�؆�S>��"��B�G����J��hNkN%�>h��R���I�Lؘt�,!H��W �h�V���:"�`�6���N-��?36�k�+��q�U)A��K��sØI%KS�d\n��G����*LK�.C�'"}�[���%�������r�=�6��0���v�NB��QL�ꛟ�<.�7\�����6>y����y��,P�Q�I�r0��$�1>qؗ����_�%�nJb������	�����	C�H�/@�nx
K����1ѥ�k��]���@��P���?��"61�iU&\�V���y7@������Ǭ�2b�x/�w��j��A���O�<DO"XW~��*���0'�`Y��T�/���h�g	"ZfOA�E���� c7]�4�<��?lRM�Re�>��(�]��Re�����Z�	B�]��
�9O�/��D���k_w�x:�y�4�{C/��i�M8I��Wc�";��]�dN��Id�e�'��8vEpK������G�����L� �:�s
��k~��!��Hj��:������`:ő0�6XG��`l�Ժ�LhHˆ\(}�l��Y�+I4�=�|p��xz Y8�����63�Dn'#��
Zh�������*�-K"'���A�Ƙ���i#�.;��^��ߍM�=0eK����Zn��'!���:	6Z}+1FUn�jk�%.!�j�}�ţ���Ky��'����rS^��%�tT=�h,%���~eh)cO�	�|(��7��ˋ��F����+��º�*�{�3`$�(6]�&Qi�+�m���d��%\%��+~����4˙�#��d�r6�:yŤN�lp�!��(a0I0VEp���(�Ƴ���P&x�OZ��{�9�*�_#һ�#($g���u4���)�͚�&sF+����x#<Q�P�7��g�����,=H,��a�ӡ���7	�8�NF��$� ��c>H�,)�c����IX��cI?���U0�X*�������Cly��凿�m'�+5�����h��L7o_�����n?�t���40VҌs�ph�9Q��%���!EVv�4Ex�>D=jh��/��o�r���;����fcR)]?:��`:*j~������R���q!�;&��J��6����K�R�-�%��!(B��b�a��P{R���n������fH�����+�6q]_��?�'�Ϲיt��K���H׀����n�ڢ#�M�9�E���}ط���N�d�-������*ԛ�Q?T����m{�5`Jʘ��L�iZ�1�[mn�Q���p7�߈���L\�	L�Y]�!2���"��;r*\�CG�2���d,S��#Kp ��Q���k�k1̇rH|֪�pЂ�Sa�[���*^��<�."c��H���5���V[>���Ǎ��=elX��Be&����la! ��\��U>b:���74��{YF4�n�v��4<BNg�<
M���h�s�aj) F?�4H<·]�>�M����;A)�77�$a��⩶��S���ٔh�`[d�s���"M��EN������'�B�8��&��o�n��׊��6U4��j�o�4�m���ud���/�`���Ĵ�b׳�:r�dg�T�6z'.�Wㄊ�|�E�wd
F^�,�����66�]n�yG;���Z)�	P r��_ä��np}��,,�YS���T*o��6]�<��
w����~H��3��Y���?��E.�p����8�}�.g�/�t���BJ``G���30J�3�5�At�ȭ�Y��a�Y��x�.9�-��X�4ZM���w[��9�&�f=	
�\̋d��@S�p7fƦ&;} �`y[��슋^�Gg���sL��lw���M5��Lw�ɼ
ך��k9ls��(�J����Q.	�!�:lw����h?���=��R�M2�Vp���#��V&���Ȅ���;#�=�W&`�3\a]�a,-���<�^�6zs����I�jzz����TM��#�9l/c55h�Fd\e>vY+���ǒ��s.C�dv ��Z6��Rm�5�Ř�y�'_�-��'�]��ދ��
�`��2�M��_n5��m�X���~�`u��8b����w�� 0S��EK���@*zG��&�8TJ���B����wo��:�W8*v�[�A՚���Y�%�!M���� I�`D&�m4�ɒ�SΙ����Bj��N:!�}��Δ�6H�^9�(�&������a�1�jg7�Ύ�Eǣ����t�=�^��T�'�~�G���H{g�(��/�?�� \D���p����IQ�y��^�G!ΟMQ���ߜǆj�����0�S���e�p$�Q~��mx��� Q.ncX������A��b��ג+K����p��d+�U�,?)LWs�.O�w|�b���$V9���[��{@��n��m6�ѱ�oQD0�]�1-K�)��Ŵ	4T!�T�cK���4�YDU�
����U��o.�ڏ�j}ZrtO�N�|�ͱip�'��Ĝ���ʱ�^ͥ\�HE��3ho?0~S�q��������=+���X�|�Ong3�.��o�S�KJ���Wt����=:�0�Ҧ�V�n��Q��S�l{���T����Y	�D�y���"c��b���6��;���8���Wwp�<��W��[��"i�"9��QE�A�z�+�J�����X���3�۶\�֫i�����&�d��Vqe��Dx](��B]�o\�Zuiҙ���!��'r��rc^�Ƀ���)�-sQ�	\�ӸI�,f����׈�u���3l��1���A��x���eL�m�{f�hB�><�"Je�����j�|�8��$�p�z.ly����ˏ�e"�P�O�h:ퟺ����d�}�\m�ʆ48-��*\�)raLL6,����ij�C���hI�)��r�G�ؽ�5�P�(��1D�:�!\����ʕZb��~��Ňf(�J^��j���Pw�%��)~w�����jxA��,�1���+O�pz�8�	�B(^L���̉����Z?��KQ�/�� ��S������JԱ��Mg �"�8�IH��%�抩�!��-G`R�>�<G$�������)�r˭.�.:Ee�$��n7Yq�Ȋb0���]��^��5��[?��Á��l�j�{�l���w�cN�+t�_P�?<��D6H�uÍ&ο�Ww��ja߀v0R��IB2�K��5C�7+;�v:	��T�ց�����Isc���`|�x�� ��p�����P���a-_z�����c��lc�f�6X��Vg�#S�Z6�\��l/G�[��H{X�����q:e)g�C褈a�2�z��\?Vf���,��r��LdP\��s�s�w�r��l�f���XȤ�������ԇ,��h�Ib�;cT�v�B�5�-��vcp�
�S,O�İ>�}�tgI(�=)��~�8Z���Y�GD��T��b���Z����w}�����0�*�vv��'4��9�0�1૥ə�_���n���t�doIަ����>�'���9a6��F5��;�2WC�55��Pt�i�~K<�FhwC�~H�\��f���*+µ�P�g j̀�g�����L^�\\t��Ͳ���#��$�D	\{0���ɔɒ.�g�r���
�SK�#��,F%��sO~��V�cnFM=�ǧ�?)����9w����>�+��⫺Az�郴��Y�k�ɒDG'_�m�85�ׯ2r 1J/�MƘą�Ox�
 �z``�hG��Q�(�2��o 7Aŧ?��ҙ��ref;����b��/��ԑ2r^D�3������~�w�KޤbL��J�1L	Gת�A�rdK��L���9D�՛�>N�"Xנ#�Znp�&J|E�z_p�7.0�YFe\��t���l9�ǜ�'d���
3
��������s�>�p˾J6��������M�|8�SS��u|����+��!��n�n���2U}_�Wv��a�!�v�\�N7�������1��Z(i��[gMi����h4��f<K��絾�y�|8�B!%�B_<(r"�L.�'Dz�d��b-�n�|Q�q�r!-�O��z�K(��I�yT�Å�V�Xn:�}}X����������̡����#]T���E���1�`0Ӹ͘�����uYC�G�	�l�+w�����S���g��e¢=>�zi,���S���Hvﺈ-�m\<��r��0�V���J'B���	nz.�l���gٶ�K���6%T�َ�!��� �ƞŉK ��d����^Q"݀�,�g�r�+J�z���Nz������5S5�����@�Veq��J�B����=�m#:�����,ݤ��
�����x��w���O���|lq����7~�3y�e�+���T��񆡋��o��;�tA�_�%���N�W�����v��yE(Z
(r2�k�O�k_��]Q�/M�)���2Z�fK^{gK���M��4���y��w�"�I6�0���:��D��8W���U�;C܂�.�MC���Dca�'~ħC��w#]�D�Z�E8Tە�X�~q$^��p�Z��n��Y@���^`�sf�ѓ���`]��h�h������ZT����~�;\��wʌu�����(�iM �����4M��2z>�[*��&��t��z)�ك�69�-����sG��|gy�>}	����MAL���J��'%��^3K?��q�UZZq� �fT����I��G�`I$�j��(I��k���!� w�M���ؔ��1 M�sp� G�柨]Z砺d rښ3>�HL�zב5'o�/�u\Jh�(o9�͊4�&�U�u��h*�1�I��ΰ��UpE���`�tQ�0�Q4�:��]���Ĉ,*���Zu���MR�)���$��E��.7���-46�R �v����cr��<����l�Iq@��\�!��s>Ϥ0(�L������iڗi#@}�M�Rѭ��3E:�/Fה$<�!_�*;}ļ�S����o��K�����*@
hdZ�ꤍ�?/����>_���K�ˬ#_fq���,�η,y�摛����d������O	���Bv�S����MT�����n��d<�z�?#��B`8�rZU������Qߙ��Y���+,b�d�9j%���ѹ�U��_Gn[������&X�ᴻK��
c�'׹��!u���H��%	�j�nl��ˆuNl� �ZY����=3�w>O=��-	⃴�~P��y�qMrf%R��^�����a�H����D��W�o8��O����I�᭠�K��˘�aڱ5+����5�t/_4W����m�H=�ՠk��������n���Q���tNG�]*�
\���8!Pu0M\I5�<��9��l���fJ�lL眂��M�U�Ӗ��+I��/�6�5t���򭨓q�S}4���óY�H1�02"#�P\�\<�����1�\�1
�"{:G�F���w�<������,�ei�3����@1���0�J\b!In�A4�á��A͛`1_�����Cf�Jm43�c��c�n�z�@� �T���E�2��6H~d�Mw �C�jl�^�:�����۹q�V/&��^�|r��{��☽��UW"Y���"W�����o2�?�b� ��	��fv�?��}�?�&��ߥy��
�i�&ͺ^}��d�VƼ�	����83"�GL$Z�(,�G�P�(��-3^1�˔�����wqS�
��w��k�/4��n2He�/��L�A	=���q�4-�&�?�@=�̚��jv�vj�V/�����¿�U�&mL�>`3��*q7�R2g�|x�.K�Ĭ�w4ۯZ9;<����Q�c\�>aX������UQ�`����1�Q��e�j���v���S,ա��D�ZgA� y��ynL�$��6P���>��;Jj'�|�����zK�[!�*_H�ps���1UL�f��xD �_�y-�Z�r�UI"�9"וY:����G"�6���A`���ėw[�x�B]����p맣m�{��i�1y���D綗����(����l���ڊ�y���&ɧrܭ~{|��s	�*>��_��m����`k!h{7�W�$���@�z(`�4��7�M�.bI������̪9r~�J�����!�@cK��]:��)׿������&
j^���:PTV��{�d`�$c���cT��z6���ݻQ2t�3�*1�)��o��F<~��\fh�����*���Jma�D!�O(��s#�!���TH@HR֜N+}rfD,���8�a.WH!�O��q���F����Z^��B19kz�#��ӧT�G�s���vK�g=	��\^Bے�LFd�SʓF�$rR�ά�U	��1=�wl�M��+�sV��i4�ʝ��)��&�;m��-̀�Ϡ��Q���'�c�y��A��ʳ�=��n��5����E_���c(@�S
+�n�p[#�/�2�ʶ�I}O�e�|8C�x�
y���P?�1@�~=��)z
�Q�iU���fgu:8�%q
���� k�1'�8��\�@B�4����n�2���l�����˭_m=�n^30pٽ�,ѵJ5��=%�LMU��rh�����Ұ����A�ڥ.����)mlv�k���59C�AZ�����ʳ���!-�AyҨbRB<��{��h�M[ҶK�p-�[<[:?S�A��3vع���"A1����� �������-�_M��W7&I�_L׎IY��ۢ���n�N�)���ޔ^�K�怮�U�1�ݳ�nU�HE����R��8�0�>�M����Z~	� ~��%�|����&��8�3�n	ݭ���8�,�-��L�%�v��k����RA�ӫC���kQ�>ɵ�z��S(&�X���\��#�Fa�З����rP��y�y}y4�
��Ҹ�n7<`:����Ǧg��"eK�U�a�����h[ǀzK��}�\Ϣ����<X��$(�<�i��2�lV��/=��0MR���SAl��a��[����]����׼9��j?n���B�@��=7pW�H�*�>z0���SU�#�?�@��G3w#<�$Q������΀�~bM|8˶�՚4���;�J��#��(&0��w�@9>2B���s� 
>�\��\3�F��,��2k7k�l,����w?��� ���o�q�j��9�Rf����'8P�d�u�f��*���'"5����m�<�(CR��7��[��������|�������Ȁ���kFo�����y.��Ӂ�����'�/��g&�S�_�ԬJ�+)�g@�i7PΑ�����h2�G���(��?a��hMm��*6�lvh�h���jJ������4���U�憶��[I�Z���&����*�gG,�i�/�>Z�K-M>��4�jko��s�!�=��[�����Et#��2N��Z������}l���U�St
��td�û��1��<�7�2Ǖ7��"�*�jR.W�R$q�%�"-^f	�Nm~K�k*���M��L�y(OE��$e�:Q(��"�Ȯ۾�P����Rn3�ִ^ݰ�����IE�8v�m=5�lCB�e>�^{�XXi%oJ��ۇe�oo�=/QDۈ�a<&��it��A����Wkm �v�����|2)�|-�<j��a�B&q�Oz
c����.%vQ���b>�NB���(R��o��E؏Q�v+_��퍟�J��
�U]�څ �E�7��涨�׊���(��䔑j���%�x����h�i)~ҿ�L\����4�wM*�Eb=e����q��}�37�uIUo�9�v�PFR�����2+�:&����P5�2��R��Y:&���U�ۓ8t/`���r�j���ґ�Y'V��ήF��:j���i��굜bvUʋw?�v�)ޘ%G�L���돽r�̪H�k����v"�/�;���{�:�܀�#��?���')���Y�9Y����������`��v�,O8�8��3��H�h���ν���m�7;^�5��;Q��� ŦG�ƊRU�f�\�T����}�Bxx$�xS�&U!\� �<�F�?��{�[��3�(Z��Ǚ���a�};�I�zIh�9S����(G�/UF��a4�+��v�Ż`�%����{�',�������K����9�<a�[�#(�x
���Y��
�C&���O��Q���"� ����Fٺ�:reP(kÑP-��t�pu�k ���,N$�8��E�A4��Xe�6L�-�d��ۉ�UH?0���6xy\
|ŧh�i��{���f�����|:#��eQq�����:
��ٛU"�%
H�~�p3 ��;��I�T��/�a��1�=>�p�}!�����#���c�:��U`�00#�;�5ਔ~H�"�JY�E�z�L��o�*���1@����Ӷ��М_0���ЫÖ JH���Ӳ�nt2�C�qL�X[�e'��Y��ĉ\��	ћ��;�Y��_�3�z�fHܮ<�Ͻ���S�5x�L3�ׂS�Ѯ?���j��υ�r>9-ğ��ur�z����J؀�=�7�v6i������-.�އʊ
���(	Nq�x@�n+��x���L����ޘ|Mbs:��3��p�� �:��7P�s����U)�b�|6��ޒ]3�oz"��f[.4ϔ&�"S�~$������B�~X�t5>c5�N+�h%�`T�x ����Z��HW��X^4�[U����
^'?�2pt!%3vnN�j���y�e��b�JP��) ���%��ڕ��P�d�Ǿ_8���yhZT�x�D�B��M|?ʴ����:Ar/<v/	�V$[���棳D8�P �������q�Z��z�8�9�����n`���P�&e]��E��8�
v�jU9)Lx;�7o>m#i����V��� S"��|�Jv��ܿ�7ƱM���B��\�V�]I* ���0��%a
��2~���\/�&$��x��2�
�Է��D1���Ln��{ܐ�J� eVL���z|pQ�;���D�,���E
����=�%5]�m�������� ad �}�Xn�����&��n��ɣH��7�4��c��13MIG6V6���8 s�������[�����KOů��h�6�#�%����z��5MY("�����c-ALD�����g�w�s)q'����>�vf�W��A
��߿ohb���E3�	=�t٦#�Uv2�&�N��I{�hoQ�k�xm|��{��;�@�����H����6�?0��q��Ub�ee�N�+B����ܳ��:{����2�B���σ��~u��mq�c��:b�	�Q�KcMe�-�j��'���z�I���K�}��i���`�V�[ F�+�\��2(��7?]cC̨$��杷���<�Go����.�a6�#�hCJ��v" ܾ3W���`�wM�J����2�/y�0$�n�(���R �5]'�q,ӊՒY��}�����W�GQ��E"\�k�V^*B���!G>�G���֭�n;S�4 *�_���2x�k����I������u�-�n7�5�*ޭ��7���8�v���x�Ux*˒F~�/�o��P����9���`�%#ߺ��{�=���N��!ix�%�(�&�棧�Xў�T��ǲU'�%�
V��jPr�E�ɮ�IL�ip�퉈�9,*�´��#���K��Tg�N�Ƽ�-����Tƾ=�;1����X$|�����ˬaR�̪�m�+L�[q��@�E�|��l�IZ��ߊ��:4]�����E`���4+�i./w0��+&��t6:�i
9�*�i�Ɲ~�-���^3YW�|*^,���ɧ�Vd(S�'s�E�f�?��nY����@@�g0�L��!Ϊ�1Y�t[tMLgo'�*�1����w�¼U	?q��?>d��=������%g|д���g!��u��Ӑu���`����
i��5�Bܦ�f[& 6��F���E^?����3g5θ0�3S���)�N^���/�vܱ�
y˭�`�δ��IWs�������ߺn�[��^�c�3;�ӯL�z/J�ytdo�4A^��<gR}�Qt<j��'��|N�Z�b �X>�P~3z�^9n����Y�{[�& ��'� [�`�4�B�?�,Cr����Ŋ4խ���A�1e�p=
����KoH୊�p1�W�0'v�(q�]&+u�%�z�P,�P���>5E��T�1�	�W{<�V���n�yM����̾=��HD������-�~��n�%�^��FW��m �����bNV���t:��
w侙�E�`�	�v�2����Թ�93=ɑi��BØέ��@�m[Xt,�]�[��ˊ���`i�>&9��+�Y롙��Ǣ�R�?�e�	[ ��B5�/Y��slY���N3R�a9���9��!�0�b�K�B�o�� �s��΀�_Tߍ[�KӖ�1��N���i.�W��l���.�Zy��W�DO7�ѷH�ܫ*g�d9��,3��5r�� 	�{}�/��A���bb�?~�>I��?����q��Z.� ��u�8�IM�=��Qt�hEr���$�U�:��� <����O�͂<����h��8y�G�c�C>(��0S����q�O�i�+m���-��܁�$$�f7�V�5�x��w��5͓@�P/eD��������}�"�����%M�k��S�7�0��룪����K}jZࡽd�i^��Q�QQ��J y9/�[�펧��Ȣb$"VS�i(�'{�^��P��=�Cy�n$�4��;����*�l�I��P��tN��O.�Dci�K]7�i�H���s	~ #�s��Ǧ��I\���|�h\t���‬�e�w��T�!��36FEg��(�Q�h�5��H�S���%�)��3�lb����ѹ����r���-�G�x��̯hw��y����G(ʍ�GZ���k]U��� c((���ѻu����V�>HYI"��8�\OQ�P��~:���`�iz~pK�.	���s�M�M�ui���-H���������FŅ9jݪ�X`?`/!�o�͵_����s@��J�a6(�Fcڹ�O(G?�8�^�@��"�)�8���!;	�GU�&{1�������)<H�Uu�Zr���e�m�-|�ئ���nk���19W�lq�-j�e~w���'��ދ�r��m�c�zjr�Ы֘�zc�z��'�wES������]�)��3�@Ijd�Jsi|ݏ��r�)Fc�������W�<�ow ]AKp�9_Y�^�P	���=�r/̸L���z��>N�p��J9�FU�ȓ�=U13�����@�F�JK
���gu9�\�/B���]K'�Iv�;��[��d<�2���8Pc6?���}�ChO�S�Y�]ށ]�D�ʪ�7�2
,�ڑ:��8?�^�������h��A����A�!���f��.�+��R�	O��v���ztm�F��)l���WB��8¿�K�X{��fSs2\䲴�%ĸO�<�a��"p�-mmL@�V����{������I0�ԭ_N1�)�ӧ)���3��ޜ	��+Y�Xg���A�t":�o�L�4��s���9]Q�h����m]{-u�	4�#��X=O���ߑ�24���9 e��1����
yR-VW]��i\S�y��sy0��C�cW���myM�
�ذ�����[ƶ����C�rd/�Ź�vw��&�5ܹ����������TsĎ�i�v��:+͸�ԝ1�B�.:���hH�b�ʶ��k�o���DѦ���*Kd���Ә=�Q���'cg��o4���(�	�]�z\�� ��Of�;x����$�1�8ۤ�N�iӺ�9I�x��:X[��#`q�X�hX!q ��ˏP�"�i�f��u�92nVH���\�t������=���&0���'275��}gi��^��������I Y���qmrv�!�T���^�����0�
��e��
�X�V�,P��~�o�:�S5����5�aZ ��e���c)�y����܈��G�US�B�]&7�tĒ���a�R��d`D��Ãl9�#�`{�r&�#�^pLѭ�.�`?��@m�@Z��>��nO�a����6W��YY�CبƨӀ����yN��, �YU�C���2�>YOu�hD�:9���zeJ&"L����zKE�1�5��?B]�q�$��
?.��;r*݀Z�É5*"qks��d�12��(���XK�$�d����Nf������x�	/Ca{Az����d���Nud8����GG�
W�@��Y����Q�iuB���ȏ"��!��=�#wFrJd��-�Ik��Z��{\����B������<����-W�p>��`
E%�i�4���i:cK@��*X�xc���0m:ZD��6�g*c����Ԡ��[|�K�Yq�>Q[�=��������3�4"U檃���F����T��ْ]Cح�F��byk��8�C�u~n�$U�XS<�ܫצA�Kz���6�5O��t38���=�(P ��P:
���v��Zm��`�Rܽ�xP -�|w0���O�*�T�P��p�'J��|K^E8��fGzk(�����tRV(+�מ��tQ��8P���ƣ��A�7g��Lxt�s!��:Q��=� ���y,����c�@����F�Z��Ê��%�#gץ!�b�c��N�O({���2F�����p�Ycs�mA��u�J�i-�<Q�`����l}n�k���:G�G7�UM����FZ�5��KxX肏�
O��i�i�ϸ��\v�x���ci��J��R�`�φ!Ӧ֦�M}_y�캤i-g�>X������"V�Ȋ��!��N�g$��΀�]6�dmϦo5c�q�mހ@)�:��Ő�5H�{K�q�e��׉�_��5U �ew���ú�0��7�a ���R���{��d�9�[���C����K� fO[���*��)A����U��$��K͝��C�9��>ƾ��ႋo�3Yl�RE�t����;_��B�%疎|����_�]�7�Éq5��m��-�����-�f�A*����N&Ѫ���)\���y����<B(?��ȯ��e�i����t���2B��	�G��Y�p�����7�`���5I��[�A|��pe�
|u�~�p(���_O&`���\�aqV���=i��A�@��K}}կ����wS�܆1�?��Qػ��ȏ��v������ޔײ�j�j�J���i^�іq�&-�xU�H4�A���N��?�:@#�޼CZ_��z���u�N�lCJ��0���X\�P��=�c���]if=��r+���~��pO���_مGy$;����2����AV�R�a"���wb�K��5M�T���Hϐ�ٖ`U��Wy�g`I�i%ٷ�ڠ.�j?帑^o����SG���Y�����h��$}�{j�$��̕{ 't���Ҵc��z6�Iw�ʟ�����EW;�z2ڵ�g.�e�_ʭ&�GU��E�ua(g�3v��E��y�<�(���� 8K�Z�D��L�/���T߳M*�߈G@s5��n�� /���B��;�N��3e$0�l��\�s� uU16f�7Osi�W3��d=
+�Bl���A	C�W�"�#�`���N9���|-h|nW�C���d2���/<S�˄$a�Idɢ[���+��pk#�z-��˺����/�+�l>�җչ�-�mN���!n���+s�X��캤Iqƹ���Pi0��:�M�_b"�����W6Zʍo0�y^���$���d�R��jo�K�¦�(Bj�-<BN���K8�A��wr8a��s���Cq� �oz��P�Ѧ�">�U�hf7ik>7^w�[rxL�>ה;���Nrġ�|�K
IU^��̵�V0[�'��W�%ίp�r���U���_m��3���n�4;��f
����H,�jկ�{-�ҍs�/��&<��ܞc҉F�Ph���'����]֕��a18�A�M`������-�������OQV��R}�m���	��Mz����f��@TJ�KIǚ��-*v�ʀ~3� hm��m����+�����t$���و�3���X�+w��~i�UL�G�b��

4����-��*�x8��_�R��k�n�bi�*iQVZ�8�K���&����mH%<ሃ�c�5JL�Z����\ƴ?���y�.��G�7 ��ȗs_��a��%b�$#7��6 
�lD�1�A��nW'JG�*׌���:�ǨU����¯�����8X@�)t��;��i����,�r�|\Qi�o�XЙ���K��c �U'aG��,ƾ�&��.��������a���R�S��3$d��9��H�$��#Le?Ig��u��_S��}�O ���_���Yo�f�*N���m2���+��;&�#`+K8�k�g&ʜ��#qF�ZNKB�� ��^�)3b�]�O���~��&+�,$I`�`�Z+)�����e	<@b����1�~cP�����O�cU�C���)�I�'gl�hm���c�S�n� �2a�û���{'��9��QT(����;��w�%-q���GdKz@�$�x�k��W��-$��ޚ0��jn����ŭmzDG�9\�dR��U�/��J(�4*�]��p��[G`�1˩��hKf����+��9���VD^޵&W�3%��/"&�y1�nƶ�ܟ��m�)��`�3�S����R�@���q����`8v�<��g�	-f}��Gv�<%�����4t��q�1NJ�k>s�g���)�Ӯ��ߣ�R�K��'�곀�%ŀb�L����i��t�A�C���p��ĵ�lp$qX�dB�pp�z6���G�WB���S�i��+�Fo9�`B0X��*pAՃMF��ߊ,�^C"����腒!ʻ瀋d�Ia�aS�,�d�(WMMp0�,Y���)�i � �Z#w����p�Ӂ��dR֦���LM|.���ʂ>�>��Ϗ�}�d؊��΋�bW~���HF��{��TK��
6ySH�KTeDB�@� �B�sc�HW8����0)ij��^�w�Hz����w�NSXq�jgy%cRTkdG�ͮ06D�j%ϩ'�O�j�@L��Ǥ�%��z���`�?0�6���l)��lµH��>l}؄�y��bP�=�K_Up�� �$��[9�נZ1u�]��IS�:Y�1�{8�������)���m��|��Rƛ[9u�ʆ�l�S�=7(��1�E�$�:w!����;�c�'���<��{ߣ�_�:�9�r}�P撷�(}��P�6��Vh�$���s��M��M�K%*GJ�=;��Ba����O����/@U����Tf�^"� |�^H@e|B4Y>�:�"���	��q����T��_#���	p����GE��pr�I�]��d
ȳ�eWɋ��K�i�6-�!�'�s�	a�������F^A�ލ�Nì33��h�2J"uƍ�H�I�F?	k�<������J���v��a κ �c��NXݵ�m�I������p��9���q�яrV+\��W���$�s}��4��fݻ%��(l?,�K�bI�	Ѳb�TQm�r���စh�\���0-D-7��RV�q2䅗�ޚ
t�b�4��pBZ��~��;��.�Iu�Qq���-��N��~��0C�����1�c�w�+]��gCCC�蓸?��z�1IUT��޵*&'��q�=�!wV�7��K)+�,�ȓF6����X�u%��?k}P����t�"�E�˟�׍�#NY/l�O2�j���r��s�)��X��S������*n����@~��&�uyX5F���ѮJ��}�<�m��n���݀���SB["�DT��q���xQl���T�8R�`��*��S��#t���ԆW$�drx4c=��'<�1���z�����X~�����CK%t_{*_���NҔ>飙���n���~�I����$Wc��rw�ws�a��ɛӴ`dۊ%'�ǉ� B�� �L�����o��с^��$�4�����u�NS#ͷ?]Jg�؂��������^��Cؐ�~�s������.���{���B|H�����49� ���uW�_�V�S�N�?���]�;.��R�oΡ0��@�v�Txp��| ͊�J�m��K��7:�8�6]F�On1WTv\�Cj�]&b47��R�Ct�?�Pw)4{J$��C�=�o�(�����L��`2,r!��y�-�~�QO�g5�o�K�=�Cx������ag�%Y���s�{��KIo]��e\�B�����%�̓}d� @�R�lb�p���0C��ϥ�S���vV)�h^����쉯"X�"�7YW�&;e_Ջ�4�t�" 	z
�(9澓�1 ��*��(Խ��	
8Ӄ���T�sgr���x�,J>���u��)�H���m7x�t��wPmJ����h���� ��q�0��O7M/W^.�c��w�帗�����QK�	�#$�
�q��6�ɣ�6e�^��2e���J��O�LJ�F2�8�	䮘�7XR�1��G�z�s�����H�5���g��u3+�bD��xb0�/�ÇInglA,ƭo(�4�ͣ#]�aZkJ��h�4 �?K̬V_/^��of<��w���M��5K�D���Pt��P@	e6l�ł'����0b9\T^�M�;)jy�u�����O���h��X*P}��=ruN�B�p$/�gO���q��0�4�����D(�+��#{�̥8GH�4��1�O	�>*�ɹ���/\��y���yC�v�ѾZ)b3���3���g�^�  �c&SoKC�=���Q��t/�7�g[�;�Ǒ�:-�6��Rw�[o�&�dA�4�5�̶��:评�SK�G�{�@}Ǝ�������I��s70�mJ�%���O�����!�#��_ӀԊA�@��w�p��~}�W����
�9��½�P�\��H�(E�a�%�!�T�[˛)H4��y7����w�K�aj���y[ޫ�=Dxb�hw�<aT��,���GGY�n��8�t=BLb��3f�8���-X���ԧV�Ǔ��S\�T���'�0�ݾ���\n�##��3�5ЊcID�D�x�^��B7���X2�z�t
N��Ҁ��zi���Td#��>� ՏG�^藾�r� �@n�.T�(f�1��O�Z?���OǼ��\@}U���nҰ�L��n.���IX<�KT��a}n���k�YZ�9b���f������?��?��QR�'���6��侯�1�`:�&	*�>dڷ��H��D�"-
5�R�WS��xf�#;ڽ.�*�LD�+?�Q^���Z}Y���������.ѡ��Y7(, +/@ͥ�JQ���z?*��'���p�&��jե���j�bR`�IAz@<̡PSG�hW�XȺd�X�x���n+?"ޭ��j[dtoN�%���c�RLxV{�դh俰�J��:j�5�:acN�%�̕�F��W������b�be7�'z���\OW�Z��Y�+Of��� .�`i�o�l\�@�!��	���!|�M����o�}��Pz���"��WH���D�+R9���NpE>��4���IK�9�Ł��9�Ɨ����_H2�W��JQ
�Ƴ������|:��^=�t(�����[F�%�U�:؇���-9:�x�%9T6L�|�ؠ�n����eu0B^�)4��y�Q�Zo��#�sndwH�֣ċ�
�~#�&�`�:�N�	VDX�� �$3�$%o����q=��jGG�a�|���7��ڧ?�gs�#$�����!OK�_a��ۊ��.���a]�!�GK:'�9�!b�T��Lm�
�C�e ���rڸ���ȒW�T��*���T��2M	-t:��� �l��@49>T�+VZ�਼�r2>ƭ,.��*^�H��K|3����.���ZU�*�=��x&�o�</��Ԫ�F��5���<ޤ�Dq�%�y����n�TlF�B.fV�gd�m��?җH���_�c��L/~q�\'v��Ӡ�4���R�`����b_�bm�^?�|}SN95��n�(1g�4�������H�$e�i�x'.F�ڿ��"���C�S8�H��\%����9�#Zb��Y�*)gE��'l8��ld�r����¥�0�aKDkfAR�?0w�wsY��[߀������)��ğ�4�q�fq32���.�(��ߡ�~�"(������}Pi������?�8c#�᪫�/��	�1�.�SO�I�s���h�K'(�X��C�Q��{r-K&�+�=nao��n��3�l(��	��׭n��n�g��Tdrߑ¶ ���.�K��W���\Bý���׬�B��}���� ���D|��}��7W~�������;T��-I�C4��g1���{�r:�	S'�dz9�fu�_B�ur�X�.���,�_���2��3c���BiA��������(��ӹe-A�@w<p�/!8�0��8�~7o�JK¶�o^��z�ã��m�5}��&	�dM��<N{�}#��s~V�f1|7��wv}��;���f��Sp�[�I�|����\��)g eVn�dc32��ӵk�E/��	�����c�mL�g~{l"�����0|��mqIrx���ʙ��=���G���=ng������k�����ۥ��?�g�1
X���c��%�Kͻ�d"W4�m�x';���Hȿ��l>yG��11S
ϟ��տ�Qi�VR#����iBc_|@�RաHaCm.����ɖ=ܿ8p�c9��(#_/À�<��M�R�|���K_�����KT�ӠlFrK󠑺���(�	~.0�DvdJ���M�.��po d�~R5ގ\+��c�?_��}�F*��EB�[6^/Hc�t�|�Z^��i��$^)Iu��K'G�J�����H'6��?������kiD��<E����2p�@y���e�*��j�4l�3	MFʻ0�27�˻��ը��nt� [�HD�|��{')s�����ZՍ�oKn\��<~���n`\��|��R�:ُn��θ6��X��AZ��p�ER���V=�Xv�^}Eag�Պ�ɿ��@<���VsRbܰ�Ӂ��c�Nh��q%Fhuܡ�w��i%���3�!��#��������ME��^	��!�D�]<8Pi.��⣠S�كbD纘Uo@p�%?�}.����h'6��ʻ��CTiE�d������`������I ��E��.����T��:�������r��H:-F���3Ms��~�K�M6Ӱl.wiw1Z!X �1�L���q�����WO����%�c뭽��E��@C� fUFW"3�A���n�wƤvn�4��U�|�&�����	"�	�,��/.��]2JQ�б�ݬ���&�$��b����d�BG����)ԍ�\����ADB����"�kK�DT�"d����,�
*}�����P�TƎ��;��RstC�@r���f?�M���vE���
�6�?��_tʭ�Y���*�\!�=C�h���j�|ah���`�Ku�C�*��ʾ�Ʉ��F�[^��������&5�s�c��֖+�L�p�V��&C�&�1�s��2��y�[���-���2�J��߯�TR/�
û���CClV���X�B�խ��kH�O�s����^�!�j�c���/�g&'�j��&���ʜ��
O���d�U��a���ɗ1�#�A�gpN�D���Eq5 �\��SfK���VR��v��Z��6�N��^�OgU~��t��S��z%�S�fHT��8����Xf�&�*�~�3�[��g;+����2����<AO2�a��O�䎐��d]��7��&�h�����i�I���݆������+�A ��h(����yGwZ[���[MZ:b~���F��1ey�o�.n/�4~�E��U#(	/*os���!�Y��d���;�ֽ�̇�Sc2��|��p��5��!"-��nate���=h��AE�=	���d�����@����$��ʠ�Ǿ��a׈]7�]7Iꢀ�vS�C���V�U�"Bcl��c��lv	u3���F�����^�(Yi�L�Liن0���r���fڮ!3�v���n�R~�;.mW&�cDs��dj ���7��9XD����X�U9����Ud���r���{*��C��óH�9XS���|L�[0j>c�i%���H�Kr`˛.��g�v�	R/>ڦ���Bw%W�*��q��h���G����t}����)q��?{�",vulM�r�Vj]X�T�\��!���5�8t��:�^��͊���!|��NPD�߱���o~ ��")F�IϾ�o�3z���1������)��rp!p�/"�l_w@��)�y4��,�>�^���l�1�p]��m;{�D�nY�_1�?'v�SJ��i#�/��_T�=|��~B_#�Y^⚼I�7?�'���%j�d�h�)��<ިmC	�6a]1&�����4<�g9g���7������̟ͻ����
l��) Vp�"ڥ��i��)�.�_�m�3w�E��|�q�9�x'~=t�����ki#q?*��Xo�n'���l�M9"�lg�Ȑ'����F���iDdX�J��(��-���ң}�.Bm�1�7o_�>K>��n��ѾF��R2M��ӳT�@�`Ͽ�:��S���N��8����GRƼ1d�'u�d�{������K���+��2��A���j������7	ڃ�)Y��B�̤�/�� ��Ayero�m�ڲ$/�|�$��jʨIN�+	�Q�G���xv ��~l��J�z��t��P���-�����he��{VE-���B:�pO��#ؾ��x�;�[�$�� �"u$U�`��� 3��$���sBGF}��<�IL�9�?:�iK���t�d!m�J���[��Wi2�*#r��9��T������Dʰx�;��1��2GZ��]S��۝�<~<5��f�K�&~R ���lK%�f�h]E���>����n�6��}@�4�Օ���������@V�m�`Z/G��ʏ�G����_� kߛ_\D�/���xC���_��e����= j#�앏���ݣI�x�{x�e0�C��"�W� �y�r�*�<��}�Z�7��l.�	�<�\��t�|���u�K�m��9K��S`,m��RQ�@����K�ɩ���87���w�q�>z���q�hd�����X
�F^	�T�`��3 �k?����&�c��VѫӁ��l��\�xb���9���A��p��Y��c�"	ށ���R9�S_p�~��*j�˗���͠N�xHo���R(	)/Iu��,?0�S�E���t{�ĺ���%5�!j>Į/��j:���fM��m��[���-��YDT����H-1uuҖ�H�Qt���zk��x���ж�9�ft��=1N���T\����A�O��wk� 7Zw����϶�!�'u��b��{��|^�Z���7�alD�{;(_]�&�~�Ja��vP~�B����#@�w��j&b��o@���*�q֛�c4���T�f�$�:^���6M)����,�i��|D]�֪Y���|�Uh&	�^2j|��jgz����}E��qi!-�� � `u�W]�F��˴D�R9�VG��$^�q�v�5��f�{�1c�3�Ĕ�̡�9��a5�7яF���J%]��a�αR��
o�P�%�Y��ǩC7��M��u:ը�6�� ?ds�[���Jr�������l�v�% ߃��������ј܎�t����XOx#����	KH���H9|�0D�򜛤x���#��c�x��(\�5I)Z��zN*��m�	�cU]�8��L�1;`�լ�+8��_���G��Qz�O�A���N�G�9O�
�'S8�
���g�E�
c@���	§!s�J�m�X��2�%ma�ڿj��rLk*�zz!�p���uI/�ǽT�x #b��^)ە�'w(�ʴ�[�]���2EV1	{�KY6�z����p��;����F_W���ŕ�<ؼ�W��REC�=
]!6�f�����*r�[3-&Ɓ�g�r�"p+�",1uo�l�n@�>$����C|ON�p@
�ؾ��T�̧��7L�>.�������A�ۧ���S�
H���`�( ������I��P�D�m��ŷ.�=J1UZ+F�L��ZM1;rB�4]���7������O]C�O�&@P3����E<�
�f����8��%�״t�	��m�1����Ī�A�r�F� w�1�w���__���8v��/"c˰=�T���� ]��=Il�(Fa��EV\!uca5� �A$ ����M�SV�m�{��ىE[��^j�/H�k�3�b��8?gp��ej��G蝓��j�"z�����^ɶ�&�?��P�b��iX{�_���� nL$�/�z�e3+1�)����̱3��|2I ��Mr��u��O��#�O$WD* ��	�8�7?P�̄f��Ys�5 �χ:L������2-�3L>�N��H耔�Y�j�Y	�ʺ?�q�Q㰳ͻ�Y yV+�M��lJ%M�4�kQ�������Ry<���������"e��oBF����5��+�[-�8���R`�_�[ff[��4aD��a��:WW\�dK�7�k�k�l�_��3-�87�j����%ѝc�C�U�Ѡ^��L���8&�v�q�NM�2�]�}���9�SK�t�[�ݫ�Wd<9y��m痝��	Ag���ύ��w���V�0k�DmU@N��L��Y��� ����t4ee�QW�T�������C���Ќ� nP~�*Q��8ٝ��k�:��1�T�=fz��Tor����+�q�b���3������w�4�ŭ!�U\4JoSoA�!iȍ�N�=]��ּlչ����W��w�l/5et-+P��>ў)��Zdc>Ÿp�ti~��e�~�Fi�bK^�=�}�BO#Iۑ���0�d@��2A�����w}�z��)VDe�8Ji-(RO����1�1�<p��!�]F�rә8��ݚ�8U-�WO��m�wU����s#/�'b�r`+�s�O�{dv���)"y����eǒ������epz�>�2s�3%�ƲcQ���Si��#ķ�9��T��?Ŗ�
����1��À�KMC�?
�CoY����)x-��%�2;5��0�G��7��* �͟��!�l�p�Y��Ȯ��6KV�PM��|N��U-��Q,�[�En�W�}�,��ׇ�ܗ�r���m!��Iǀ�E�E	�ǐ&��<bH����q�f��� �k;�X�7�4�(J��}�/�i�(J�&���f��kN���%Aɕ�Q�����d��7���V=l�8,��U.����Dx>���,�3�k��}�f�&֛'a88|?�N�%�!2��l����/S6}���G��50�ٜ�ɇ�E7a���Ϙ�or�5ˤ��n�ҟ#ؠ����OF������a��|H���t5�YmG��K>n7�g�k�S:�ߙ+��/m�x)�ZD8�o$�w����8���O�G�{�RTSA���T������a�-R�p��U�>�/�V z�n�7�$�d9٢���mݧ�e�=�)�k�7`_��}�5�̈́�����ә:�鉩�	�@v��A&�����1i���}��*Ҡ�(,q5k�Y*Q�N���ELĹ߸t��ִ�e��c���8��xſg^�l���ǶC�����J�g�f$�Hu�73qm4	aO
�D�0�wZ8-����9m�/���21�+g��*�Ig�4$X���H ��6��Z��Ӛ��V��s���޵�\�+�υ�wy�T;��G��2WK�p��>�,H�L�I�>�X*c&��_�"�Xqc��R�,����&</�	�N�g��3�� ͈�{}�] �@?5�3��꘤��_���L=���>S��~�qQ��]����}�J����
Ԧ�Z5�Ŷ�C����Q
l5��*�Gǻ5%�W-�++1t�K��Th���r��g�Y�ǉܱ}p0.mBYc�\Ad6�@�$�v7p�� ����=��o�D����}��y	`�����s�<�m�{�{�8x?h/�Q���Y�l����8������`K����C�9�4]|C��g�;�l����j��&��=n�Q�&Fg�e�fC�(m8u�-[�P�N`H�5{�:{���v�~e���A�nJ4On�`%-�(j�궶�>�	����y���XD[ޢ���n�:�i�h�z"�q����9P���4��{!���Rv ����Q��鶫+,z��d�����tZŮ��:{04�ɓ'������|c��!��r'�Q�ha�f	wQ�k��� SNT�̴�_؊���?6�}��b�=C�S����r����`Q����p�ǫ�lh��^�R?���O���𠖪�KwVs�V �b�Dt}k�$�L�� 
h��| U�$���^���s��$&� %�0�ߗ�L'��ݟ%N{�>!h
}�[�}H�!o�0I�-��p,VS����fi�r�-����ݡ��K ]�g�+�A �r�)���j߱����R�~��Ul�����?9
?0ݬ�wG�>B�_jP�����\�M��A�z�`P��*�q�gET��=!��.�ϧ���	[��%�r{�����+ ��t���=L٪�+g'?��=����IT�5CI�����=���T�y�"=X�# P����-�qv��?3�@D��W0�bQX���&)ZH���E61��F�ɻNz�z��(�@GR]�H����}>7�E��5 f����2F���YL,|�����4R:EMFo��h2XLFW9Ř�w��2�+W��`}�F�!�r���y�4�݅��Mi"D�b�}���_�<��nEgwՑX<�[�n]!%e[��B0��B4��v��N*��3	�Lѕ�l�޶x~��۔k3�\�B��,��ã-����p_ϸ�w�@Q��h䶡A7+O�dH/�6,��n �VB�w���B�C�v�J�Va��gcz�E���v �J=yO_a<ȭ���1�G毊 &j|	��޴BMK\���x�?%��:f��=9K5��<ŋ%�ߥ����G��6�铝A�֕����F�JU�.������`tT�}#��� (�	j�'߆Z���5�Lf������Ã:�n�YUC�5@��Q�_W��X1��u,���\���@�M=sު�����LJ~[�<�N& �|��3����S��I�߹6�~��������+4��V����jSTݿ"!���8H�:5�)h����ƩV�T��
u���ˆ����K�w��hB0��E<��}��,ӷgz�)(�ߍ~��R4�������U����*#*23�^���}�P��]�5�Ζ�/?��M���fsJ(T�/��,�I���;,��a��߹��A�$�w�(M'��Ư�BtR��<������s7�6��qup{`\[�4���UH��G�ǿ�=�Ē�z�?8M�{�m��44�iyۄ�G����J���1�����N�5e�PQ����X(�
l���I!�&E�"�r���k�33�������7y�s�����-��m?%/�ER������Wͽ��<�":>��hr׼D]t�%3��\pf��~��OHF��N@��o�T�u��X2�����]��?Hdr���.Uj��'�I�N�x��8�$�˂Id��EV�S_T��L��Q��!`���{��&���	�%�(�u�a1,
���.�t�2{�Cy�f��ɺH��,d�T�j�PC�^>'�át��@�Z��q��ԭK3g�����$��L4��BkC��%����x�ZsnqO��a���@��P�P�ؔ^�	yV�`�G�,`���*aA{7���"�w>q=� JO\Tn�A	.�91����Q���1Au��]�6�л�����B��RpKV}U_Nվec/y$�S�_��t&9}�~���p�+���-��y�������٧DNTK2��h��s��� 8������㰐�]�vFТ�#g���즳L�|8�@��V�(1��c�� ��n��ġ���ӟ�J�*�����(��P*���r�Oj򳀖A�p�0��d���dy"Ԝ] �Eꑍ*#�S�_�'���L�j4c� SQ�����Q�]���@���X��h���PV ������7��X�0�g��1>��S�RgS� � ��lf¼,�uY&R���x�&��8�]WI��b�ֺj��7����6E�� ����J������������2�m{�UG�B�>�;���TG��2HY��H����Ǘ$f?�7z���n�g>h�4[�mH�o��I����t�i���[=�-���_�B�ۥ_ c��1!@BH� ��`Dq����I7t���+��9�ȩ�o]�p��q�i1�(�C>�쨐�8\���#R�]���i86�кc(C�$u[�S�W4&��,��YY��"�"kLw�k��8J.F��2�%D/��-�k�Q�I1Wg�)ֺ��)=v��h90Ә�𠞁?Gx�?�g$��@;�%gIQ�@��з�a���-�k����I��mć�k�?�~O�ʀa�H,v�G���!�^};h�k����&dD��J��1`��ŵ89�2�<	p���y�gF�@��;*��\�\��s)���"ȴ��~��S�Sc�K�m�4�Q��Xzʲ��=��Fq-�"I����2.(�2фC�='a���a~%p�G��q�.��al�����@�b5E�8iRpba�]Q�o���1�E����!�<��w-���3ִ%�8Q`�*�#�2�|D���K��/��=)H5�`�ea�|4�~������=�#K��.�`�~��%�z���@�\�,��$ǁK��{}��([�D��ʪ�C��r�J;��#B��-i"���ߑ9/%dk��*����%�D�T:���M��2��~����L�Q�.iվY�?�}�'��=`���|ȴ����ԟ��
�g)�3OH�X������β,u��nG$����F<��T�+{vɉC;�\��
h��.�%����9į1csVs�U�X���EUAh�u�Cw*������)��Y#�+m�17�l����Mr�@�����ovϝ���×��Np�'0�qc���Y1��ԛ�Ze��4��r;�n�]X�A�)��<���~GJ���4%$��K��\nX������I&?:,b3�7��c�W��Εׯ���$��m�M�\�����YPjE��6��$�E�3`�+�[EIg�\g�c{�!�*a$J@G��۵p��}�7��X[�VH����X+�գ�^��^���6���PJM�������r"_����D���2˱V�T�j��F*E�@��ȼ2�%�C!�x�`��O��Q�n��eĹ�S�s�u� �b�Z�g�b�/��؛���������Ȝ �2(=o넜���@l�>�ǎ����4Dиܼ�ٮB*)����;н%��wKҷ=B���ţ޻l�~���C�A�1���S
eĖ���F��ȅETB�p�d���:�J3�R� �[H�b�/�Lt|CQ³�4i�#W�J:�����'^1t���śld`�hz�M�	vИ�VkӰ2��g�n��)��+�4�wћ��;��qf��W�!N�!4�P� ��s�[ʧ>~���#J��P���N�\�0��L6݌Rg���u& ��\[��P�7�I�v(q=�Q�;)nM���b|I:Q@<�lz�:�%��/uJ���Z�Q�����!
u�"C������o���Q�J�a2F�6����C}��u�me�!�����^k����c$siw�+��+_�)ed`�ܶ��%�j�٢�`�ƺY�%0T�	)%�h�w]���e��B��lom�M"�U����=��jO�������G�LԮ*����|��=x�'�_d��1{�hF��H��	r�ʆDFCd s���N�q?�L�*��'�
��R��YaZ���O�p4�w;Q� ZA�hBv����ΉF#z�@��t�`l�ʛY���QTʎJ����i��M�SkL���0����)�|����e�:�D!�O���z�=�	b�`C�|m�N>$7�<a��q�k?�"�1V}�gmBP@�#����q��TX,pXS�m7i t��i	�1m�@b�4�
�wux��o�
SvN����t-��F��FS�|���~
Y��lK���{�p1�gR�p�5B��$����WM;���|]�;t���_R�%��\�K��0"��-g'��C�Ð���a(������q��O;[��~;�8��kQ�4��{�7u�+]�.�rZF�򁬩)�Ƭ&rq:<�|$F�p%MK�]��a8�G���͊B̹����ZH��ou����d���X
z���>>��]�Wb�J0j���i�[�¿A¢���6	-p�Ç8��+H��XXa�5'�*��#�YT�22�:;��%��Uv��,ۄ�kW���?�����Ml3p���R�h�?0/� �fU��!y�ց���X��G�,u�ёS��uSg�h�G4zzoz��[l�N�n���h+��$e�KTJ~՜���}&�6�;��6���l?�>��D��am�W@���E-U���̖'�8�t��6�,�.r�HHr����\�b�"��9����i+o�	B�k�2�,��ER��l���}���2�~)���i8��SCR��c��Lm�a��?���u��"���*#l�I=�
@���S���섻_�j@�z&;U|W��j�b�1�4���o~�I4*��x����R�R���YI�s��+�Ӱ�VR�I%�f[~b�ܚ�ִ� ���cR��hsmB����a&��|&�W{ǜ���v����r;�J����|q����$�S��Z-c�=.�y����¬b
� ��U��/��m7cB#j?��.�c�Y%�0�"��:2��WOB�'��o�#��H)�=	*j�S��2:������l/'�I�R�k�\0�:�7A�m�=�r����V��K#2��r�����u���Ae��Nմ�	zMc<V���B�@�A#;����h]���0jE-8z|3T o��3~���Եx 8W�C�3�۳�R��s�Z��?����}eʀe3A��eb�6�-�S��Y�X86 �4� ��G���2��}no��@J��!P1;t:$Y�՗R�k�L�)�� �x5+2;�ʤh�L�Pv^$�YI�<�u.
��;p,|̷��L�����zl� 8�q�f �jw����:U�(����]ꛋv1���g�<>!����h���������SZ��pأ��q�d���ޝ�1��=΄Nfߢ*qc��Gw�^��W���,v�����#�̇�6���4�|&���c^"�����Cޚ��A�xcL�zLH��{�$��Vm���%�Ky�Np��L���HޭV�=Yх����[��O��hx|Q^m1�U<E�1t����o�Uh�L`R���|m)u-2�ήK��Sɸ�O~�~�z����q~]�K����:�>@�3gO�!�[8;C�1�?6K��k1��s�� }�N�zJ�H��K��s����H�}�
��P4:d�|�vs'J{Hа��AK΍7&i�9�����0������K�ʮ���rӷ�� �>l��ޟ�������VW��GJ9�8�V�Y�$6O�`�����:Ԩ�\�����>�E�Ͱ�@j�k1ڠUr�6�&H��;�)�=�AM�x�t�)��� W��N@+��^-2@��Yr-����<�\�ݞHD=�o�N��h`CO�\�����=0�	ױ�lR�o[H ����A{��U	x/`Ŏ�@�0Vg�I�:�eԙ]����ߍh�*J#���6�Js�2j4��	U�ͪ��`B&����~չCԩZ��|&�0�H&�l:�����H
��ˆ��iv#�R��u ~���_e��s�E�1_�i"D<����I�ٚ�x#���:�y��:��4{�8h�{d)�k�&�G�S	����7�8���@�P��Z5f[��TƗ7
O8�Op�a��\�qI������We��]��1�P��}�%�tsCxYa<w�ꩁ��@M[�;ةc$K(īm��62��^l�ꩳCRJ89n���`X���|��v�2�M��8d��Z��W��)��O4�~^������V��f����F��4���(��TV�i3�ɏ{�r�I1��p�z�b��UB�^�M�u�圏*]<Nz��u�=�dm�=�h�I�^TY;����B�No*7�#+g����U��Ԥ��肿;�;ԪTu�Q�0��3d��9�� /�p�(Q���Y�2�w�Z6��S���i������㮂b��%��LŦZ���F�l>AǨ ,��9Bg�d�k{׼53�ш��Q�U���^G�r#��)�*�[�݃�����L�KZ�%'�Ɩb	:E�N�u���e�g�-E0�
��F^�5�|��
��k��7W�������Iz�g���H��o�G~Bp�͡��=}��zj��N��e����-,��8��Fw�_R4����Y�����}?R\��Pw{Q�/[�7D��?�����½LÔ���^�`�@�������L���aZLمsq�RKX���v�G>R	?l��������m����BIߎ�.��IýBZ����3��hҟ�ǌ)搵�L�9�+<м(X�E��%|O�؁̠A��=�^mPWn��F�2y0�>H%�۶iUTtj}�^�im�fj��r�h���x#W��F3��� ��	�NN#.K�Ni��f�`E�ǀY��{>�y�e�����s'()��]f�B��D.h@Ҕ��s����\?A@�/0*>��������W�+�2��!y��tzg҆KD�r+��tZQ�z�=��TMR7�)��5�����ӳb"�0����_���}�/`�J�/0+���$��������*-�=�&/�����*�Һg�J�p/?2�\r��'������ ��Eg��J
��\Lԡ�%1��d��^��\f�!=-ʟ��r��� ��@�!#�B�����3r��b�����{m<,c�/�y��1�[���I�Ct�ѾɅo� ]�p9��3�X>b��B
�.��eHP�1��▕.�	��k%c�, l�ܼşv�}o��.������ ���%X�)�=��)�к��X��Ff�&��+�����)D�5��q�>�6�}�-�JjmG��Ktc|r[����Ú�dafP!�y8��0)�\�� �2�2��O��Wf�Q� ~0)���{���D�\calWV�_��U�$��T������mrN,�Q�x��k$;=d�v��#�i�G(�Ifp�2e�ė�v�zo]�oC�ߕ���=����}�L�Q��ψ��I��(�c8��6<�/�Xm����t��dT��	bE�]| �7)6)����C`25f���@� �㧺�?*;w���R��(/����=��@�<�z_��>�������a�&��������e��Xm�ߩ��6�tc�Z6�����\�"�;s�%�J���I��-���nGTU��k����n�&%m��.qVx�����+�2I7���j�{pjʬܿ����-�E;�p��|'4	=R ���������N)v���Tco���ۉ��`�✖�G�9od�_Ԕ��^���aa�q?N!9�.(q�[�?���&_B�D�''Co(��.�_IH�ҋ03��j�����f�����,�$V���O���hA[(��I����F����I�4�H�9�a���#���:x��r�ȶ�U��M�.�X��vF�(��;X�K�`d7��0�M(��;M:}��N1��jԃ���܇��n/��쏿�c�i�/J���0��nˏ]vQ����-É�;Q�9ek��>rfN�����#�3>��T4KN���-��8�?�u��F]��6� �Ec0�)-������曨�bPc��+<��݀��p8>L.:hķ�)�_���ӣ�:�b��Bu�L�١��oŵ�8/�����A�/�E����+�UW���N�ߙ	\˰����B�s��[v��B���n�q���aX\g ��W�sF$���/����}���ȝ���"=gG`�s�x�d\A,E���(ȣ�������o�t���=%��Y��)�t�j�O-Ҟ%�?z�ǂG��Dѯp&�l$"�~��W�D���LF�W�Q?��<�QW=�'1�%$\m\�|C��|���
��q�SJp�NB	�ϲ���ܧ�XU��yX�c˨�Sx9a+��1���Kxm���~�|9�b���7E�{n��\w,�p���\���F2:�/�<���MN����m$�;��;/����S�1Wn,�d�em�9YM@����]��߶w���D�n2�N��[���9����~i��V����}﬷�4W:,��6����Q�zҍr�ą���$�� �N{��b|	���N�I�ֽI���W��퉲������%��"�,p�6O��]sʪ�9�?�(�+��v�+�L� ����U��~����G��)��F���`-3����U���i��y|��@�o�f�^Hg�4���\��m��<�w�*Vg��Χi���՟�xz�r���,�+�|��ڍoM��2u�/j0����:�Ie�7Gr�TKc2cU����tӑ<�'��(����s2!�͈�/���5�960E8	&K~�>�%���x��jq��X���.�b��P��$���2�4?ⱱ��v��,{�簞�d�C����3&��Ie�7"��i�}w9^7b�-��՝�s̬�k��u��	�Ie�Z��?��ꜜa7Ғ�/j:���IY�C�"S�)6�[K����,�MV��t�fㄌ\��xa}(�;��� ��|�:[���pRlI�Z�v�g'f�s����W�0��:��côF�b:�kX�,�4��e���y�"A���@"���A�<u]*I���oss!ے��ՇQ4�?fWp��^����&+m�L�+�um�	"��­}��vO�yW�_d�}����.���{��}.#G����1��ȩe�ڕ}h[3��g�'x��z���>��E�)7"���}/wy��F��^�$<�z'�@�e$��i�-sS\��髆A���1���F�Z�>٢Z�tj7��C�"~H
�INxyyBɟ$&/��?&V���)0^���ד�V��]oF_5�Hb ����iK��*��'��a�XN�}"V\�`��%ᠺ��'�@Ç�*�Y�]�ՊZ8K/9��Ƚ��������MUHS�:��HHw34UJe �^�-S��D�7{��5vΥ�<yo$!`;~�T^�C��@��p������8~;�����ag�^&՟���d?	~k�ĭY�FV�� ��0�n,���� ��>�}F-��
#\ĵ�RU��f�����ދ�C�$�A<�PΥ�@�XN��<��@њ��U�}�O��&��-����4"b�i���Rh�Փ`�X5��gΆX&�Do`h`^:�{�w��ȱ�䡱Ϭ=yt��Rc!C8S�*��2:��?kvXoAy���\	�!����u����*�
=()����G�,ʍw��Sۑ�%���&a24�H\��lX�)r��P�}Z�Eu#T2_a�Z8�,�w�jQ��MA��N�گr_".�º��z&��/AH#�qIl�l�����D�a�|�4�(b�|+ ��^$p>1�Y�{Ͼ�嬑HyJI*����=�fwp:� �=�_7�"@�v���!����V��|zh�ʀv��z佶e�[ɾ�⤻@��A���%C�^���+=R4`��r����Hg���F鰲;4U0 ��!ksm�������ݙ8�U�]:�%�]��-��P�~ �g���moI.6�S,pҷ[.|�@�"`ʚ�}��m9
1,g�;�̭h�z�aV��ذ�}�.�G��� �������}w��CfU�T��fq��M�;Y\�Hi__�	�������S���Pn���N�;� ���;��>'��^�u����x�;鏨�@��'"
B�aV��;��O����WGл���$]�6N���o���"2�G�恈pTQ�y��\�F��jKŨ����$�*�D�`H14�?<�錀/Ԅ���Ӊ�_:X�m��_.(S�kf-�c�sF!�	�oX�v��Fr��+�O<H���cR�**��G]�1@F{��M���Y9�u[����9��t�^_�"�3�Gv�N^5qXL�AXrӋ	9���y��%�H��
l	�����0k�<l�2Nh���E|��ҷ�����A���H0�ǎhZO�#�l�MT����aj��8y��h�>�q���F�:���C�x��*�3ZTz��`<�H(\�t��]R��M�� �((4t�_�_5yyas��fs�FH��dE�TI��o� ��R�/�N1���Fs�R�9��t�$�]*ґC�J��3<���덖��\fwsN��Z�c�,����5g^d��`��0SrqB��(�v��]�K�X߬x�����B��z��͵i�����WޢCH{�����L��:��V�_�YxYh%�:��d���^c�]�m-�?ͺqW�����5�[a����?�)�6�����4���zX亢VMsɤ:�F�~�,��Ty��"�_M�k��*��PH
�K
��Wa���tF���	ѣ�Q����,|L.G{F�����$	�NP���D�Z��6�9� ���$&� V`�I	T������,���x3��>�rm:XR�!d@eo�cbfE����;�W�uDд `h�W �+s#�*�PW�����'X/CN0�~�YN>D��Suz�0�h���UNYa>^ߣ-���ݒ�ţ�mZ{�d������	��!_%�������5?GH~�-E�M~yY��1'�P��ҧ�P���)�n:�+"��d��J��h{*�X�n��z�N��|���M_:����/�礉x֛�,������P�Ȝ��鑮eo��D�����.u&��I%g<ݟ��>�"�ߑto9e�uS��6�M���>EܽS�J#1Y7�B��L����p�7��`Dd~�Gl�`�Ch$�o#W��!\i��I�^dI�&�偼/���� 9�T�چ�e�u�f��2����8Gw�,��'�cT�d�qM5`W;�q��)AyZ�!��("���:4^��[m/�M�/��_Î���U>ͯ�a�a�B<��b֖���B��%�Hj�t٣bj���)H��꼷�4�٤��1lӯ;T冼�Et��̨!�����[�]��/쾪�F���{�Ik��L~��@�Z��֑An��>�X���c�I(�5'�DIQ4����SO�Ĭ
�i��R;,�H��6�hӭ2(#��ӎ¡�
x�lR�G�۩�H�@K�B5N=�[ʿ��C�i����`>��%HuF�2�3��[A{� ) �=�R6��iOt~��7�scY��y1�� ��ۿ�q(vA���Fq�ic!�U��p$��)<ԉo�d܆�&
/������D�% |��Z�� ܸ#yhÐ��~�w8l�3"S�^ۘ�3����bg�T`�)N����#?=�670 3�\��$3����t`:���X�\����KҞ������e��Q�(Ӡ�=�72e����|ڲ� �V�A��b�8~����~�����R�5�R�6c}��q���EZM���`;<�75�|�D�"�����I��$B�@+S��V_�8eu��nH4*���x�pÿ�ȓrV��~i�����x��xj�
d�g����u�[�v�;>��ʀsͬ��C�w���%W�� ��w��sy�U!�;�!K�P��"�X���I��W�� q�ah�?B�����-��ľڏL�r�&Z��+����q>�_o-}A�d3�Ā���Y��;��������M=e��*�\��_��RPY��=Y1�C2ߒ~Z �t�3����ʨ�'�>n�S�����jY��_���ew�F��!)#����,�C&�ꩤ�Q�8�W��*��<�r�I����<j=6��/M�r� �۟�3�8��n����.��̌��?%4\�&����I�g��r�uZ~��y�J
� 1��,������n�'���&o2~����� ���F��@����Q�~�y��FG1o��C!!���Za�A�J�Ջ�&փS��؀��J���8�]\���՜,㣍�|���=�ş�>C<𭩵��D�;Ս��`�<$7⹕	*���0�g���FX�&CQ �C���S�=�?!���_��	 v[c"ڎ�j!��RY�>H�k�ZC�ɏ89<ћ�`��<>��'��ބ�[	�1���=�j<�M�T�e��U�G6\��u;��(q�x��������j~#�+	&�t.�,�F�G�tEŒ�B./��n.*,(yR�CD����$T�vqz0�x�*mH��6G����sR�C�F ݾD�ךzx�| 2�#L��ty��vˤP��K�"pq�gc��I+����!|}%}�V���>nlvZe7�`�~�FS�@(�� nU0;
�(��C(>*�߃.��w���q����vQ��v���W�I�n8�����9ީ&�D�¯���m��c#I�\}�ӥ��vH^�����(hwM���~�Ηk?� �ߌ��d C:��X���I�&���
RaU�73�T�v�L�a��(��F�*�S�=.����[���G�A���u)��r�MUg�����(5�[M��O|V>D�/p��~��Ȁ):�!�����:N5c>gy4R��d�K�:w�T����w��y�}�I'4�8�M�9!�6�Q.�o���.��b��X/����n�)��M�E���"�Gbt}`�=${͍�촔�;�@�FF B�^�, �+�r83� ������w�~��"*��l��凯��\)���`~��zMSM��d�In���
�E���ơ�e|����J�����K�K=]���˰�k|o`�K>@
��Ac��Y^�B�.�-#�FNn��
�b�B:�r�ԆJېTP�+��2���=T�V���Ҵ��)4�Ib�М���D��j��ћS��q��	�TTQ"@�Fl����O��n�Fګ�m����1��>�p
��K����ݛ�!B�A7�|��+�޽%�Cd�-�?��-�6���w{^���O�\�X7B�T3�T[�����u#a�XL�D�-��Ԉ���p9p\t�Sf="ꈕe���Uf�jSe������,��S��0���8�譵-�^+Ą�nnW7�h�7Sn�%���k/a��_��Q�c�_�5�b���I��;P�ZOW9#C�J���_xzq�L��F��w�������pqؘ�j5ž������&A�4�q/�����o�͖���8�/Gz,�i�(`���Qi"�^廊-�3`;��g�蜓N���7t6+'b�')*�I���c�w�PH���gX�a��HfM�ۣJ'P������Z2Y��C�f�N�Eb%�W�K�(��;H��\�Pq�|�΍}`�9�)��~���Ǎ=��
�|�ԯ��iq6�v8
@R�!]ll,C��j��(�E:�2�W"���,L�V�s�'pd��r����+����3��<���N���������6�ղ @.q	�����M7\P��s0��G)V[��{�����A䋲6�2ʠ;�<�il��@1!���+���4�WZ��03X?*bX' ��-P�����B��,��U<\(�Yq�៮�I��&'�d���Å��g�{���d��z�{����������Z�~I0���,���EV)Mp�����\�g7�?��RވV1�_�{���c������P����rz�贈�3�y��7��ڈ��ǯ���w�;��/�rE���η�i����m=[_ %s���\�-�Z�;�6�8�v�4��B`q����P�*,vc�_�nH���ž��x�:���&C��l��5�N�`ׄ7�Qj�!�,��u�Z&�[��ؕ�WB��2E`�"�c��b��
Q��^�r��N$�#�,��5�����@�%H���cSK�<���cK��W�?�`��ɂ�����2f<���s�T)X?o\�۞[)��<Zx���H9�9V������ñ��'�0m��.��H��c����?�*�7��9�������3܃y�r��N�],�^R���_V<�sa���'~��}�1t�,�5��� �b\Ir&���0�g?��mu�hf�+�[�JT�2Һ���&I�b�T�5v��P�&��t%�"&�Q�]3~6���C�mB���_|dDǧ��/Y3�Kb4���= �Wd����%�(���ۈ��������f꿟m��Z똩0vW蕨�(k��ڊ;L��Qod�3e�?�"�Yt�#LP���T�:�)��v�$X����xc�����4��aa�x��?~�xTa��ݴ���h{Vd�������;5��xV���s�S��r���"Uղ�XE�e��},(G_)3u����B��~~
���(&�O��6䙪p͏>T`�[�xR�I���`,KЗw7��C%r!��Kp�!1��D���)��M�cN�LO�nV=����?��o}�í��z�epF1��,o=���5���VO�D�2��Ŵ�ڣp�PUg�V���"ı�����hC�*z���[Ys0�ÆH��\Z�'��?���/�p8�PH������ʯ�8�K����-_����	ޗ�E4z��)���6��4W46Z��,廧�A�Yɜ,T@�7��8�!�x�G����tl��gL:\N s�6��=؀��$HF�eg}�v@#��1[�U�fӵ���2M�ze/���ܯ�aÉ6��v
m���4�S�uv#�2�:"/5Ȍ#�.H��S�W�dsni�5Us*.=گ��_�b�yg^O��Q�Rm��i�}��.O[��L�ƨT�ƨC��l�]����	Ě���� 6m�Q����p�^̬I_=����~�at�!��
@`-��ޓ9W���|C���|���#�{,K ��xO"�e��X�"I��/�g���ƎG����x��A����j��3:y��W��ϣ��B�\{pEܶ�]����"��ܧ���
2�:��c���H�v��m�F���#B+l%��pfU��r���e����Y%���?1��6N�����
��*��F����5�{9�(���Sx=9[O�_��t*�Ty�2v�U'��������x��:b�ɾi��2�kޭg�!79;�*�F�'{�}�;�V[����-��6�h�j�P\��9����xow!�@+ۋ�;�mc�c����&���0�zj��iP��3Ee(�Ù��iڀ��)q:X�.:����A�č�ʹF�r�Q]��9;�/�����~� ���xjkI����Q?�~�v�&�,����v�?��%)[
�ڪ�T� -��p/]J�' 65`^f!҃����(9"rԉҥ����
��r��v��<{	��'Ǜ��d�ui�(z A]��_���H�K���
��ˆ(a�Or�ȟ�R`M��%�0^'��Bs��w����:�Iۼ��%�6*,tb�M�E�Ԁ���{���83!�
��pcU!�%�ϐ@3)7��bpQ���"�G�JB�
�z�����ZI���b����~�[k�2��̠L-��g�uYS���.%ǖ��ng���lt�2�8!Y
���=v��e���<z-n���դ�}'��ʩ'R.M�̔^&B)�Kp�P�ߜ@�`����!$T��\�I�Y�e�6i�kk'Vu�C4і�M�S��1�Ûj_݆�ɭ�@���;���BL�?�ם���ɓ�"<�|i��-�:Ag)l����Ҩ�Ä�\��"����\�xdPQ�m?����H��e��I�.��e?gu��f��o��1Ȩ��L	o�B��$�Q|�h(wQ���� ]e�,��t�.���z�����@=d}��}�~hg�ɫ�}\Pi�bɁ�::�gߜn@C�A�D�θ��AbZ�jz?&�>�Hg�nᇽ� {4P�q��,���R�RN�T��VP��S�����X0�I���Ur�.yr/�Y�����`���*ܒ*�J�B�L��p� �Z�����u�����`�M"!��c��4A�Y��B��fiVHs���[���&(�@d�>��"Δ�W�Sd5����4M���ԯ�C�cW��ep�ud�-��\ Aɑ�ď%��1�	���~(/Ǘ�-�]�,W�ǘʟE���֍���xH�1��}����;o�x!;)�\� �\��3,"�
܉)N�Q�&���z+��5�D� �V�|��ZwL���Rf��+�@@�����v{n�MN��0d��ʨ���1�!��to��g�Z-nт��Rw�uG��@��#�LXq������s%����q�ܢ�h���[�$n�N�wITSk������^��a�sʏ Ǜ>�)3��m����)�Ϗ���n]�I��-��q_w��A��L*��6�����D��H�2��ɸl��l �8�HȢ�$Ha�w���c.�h��$�'şs#�+�AoC8W9Tw��,g�G�sh������O�:��1T+˅���7���t�4`�]�k�C؋4<�����c��?߼��NN������h�^ui5��kfu�#���P�_w�&Źj����/$_T*�xt����}\�=�K�)S�=�٦q(��|�;9��@�@��C�F�0�U\�����5�<V���*��������>��V��^M�npQVFЀelxhYt$nfq�VO��#AV$˸+f�~[U?��:�����/v��k�0��F�E���e����H��d]}��W3����Sg�Ţ5*�#j�!������!��E����������쪰���(� �5��G�W�VvƬ���RK"��7�&z�&hVnjb���EN�b��F����#�rq��%N�T�%o����i܊�8��Z��p`y��/|N�� ؾ��o��]�$=*�9h[�:?��p��̽(`�K{a1����Q �h.����-�l{��ax�1%�	N�������n�*7!{=}nG�ƈU��P5e��X"���OS�!5�Z"�gd���V�a�G"����܎r�+����� "��~J�2�T��h8������%�,�Tt�0G�˦2��$@0ռv�d�*�P���H�����D��/��m�M.�|랕�z	�.=�� ���'ӫ^{���2&�X4>��i����&��P�4�g�ٲ�z�ƔW��<v��Ui��a���ҫ�^ӊ�w��c�Q9Q-��K�3'Oc�-B�~�el�["]n�0TO�
�>�q�����RlC`�\$�ԅJ1C��V�iV�M�vb�H�V>]�%Ĩ�{b�6ƻ��Sc�q0�e�*3�]�š��"�T�ˡ��w�l����gB0��I�w�׍�_ t� �;�J��/;Os:VH�+z}w&K�[9fP������Ϳ������x.�,�O�X�����!��5u���í��&���!�x`>��P�B�zͦgZ�@�X��'n~C��i*2��s�`8z�P�R,M��\��(�Һ�2-!��΄�D�OWC��w�����]�'/%�_x���<=�#�VD����X5b2rŭp O�[�а����|�*8��㷩`��d.���xIb��f���|x2�[-}#����$�,Iy�D{T������?0@N�d����\�( �O�=�E�L�J�\u��`����gA));��;�`�/h:hS��x"�M��d��H�H�KY���d��$![n*������v�P�@��.���!��!�d߻V��.���hH?h!�\�4�����b��Z9oN�z+��V]�![�I����r7c���&�RX�3� �aء���� znL�Ci���������䑥C�Rq�`jnr�zY����O�m���O��ӚeW{�n��}PoZ��h`���Ȍ���E�:MNC4)�"�yض�WZ�y�
�8㞁^G��
� c�t�:������l�Mm�L!�ğ�qw�3v�Y��;�'�� u�i�N�����;pzo�Fn��`K�;x*K�:\\z\H�u2 |�/%�z-H<� 'ģ�\�[~Dg9�[��c[�j!#z�_إ�4��gV����sD(��`ۢ���V�� J�}Dt������x�=�g{W��/tl �AMR���|�(�N��6�4Mh�aU�I��a�
�S�q��Z�D!w��e0Sc����G��2@A~
qҌ��d���B2��A_�?������eiЂ��h���ie<m�x��P0���8)��KZrv���LZ��d]E�,V$���RsY�!����>0.Yn`A e��tL)�����Q�z�Ĩ0_��1M��O8�iU(�V�4���ӭs�nx\�6#�c*��6�*_ ���W�3��,'� ����$�;��$a/�_>r�sK3-5�1� �����J"�D����B҉QR�T;9����il3�r�ͷȺ����o�ny�t��uIAGa�D�R,��l��-~��M	�	�^Z�T^g�,���� 6���@#���?���7E��u'7S����n�Xj)Ԝm��j�{G�uYvQ�5�2�o�~��UdOS����h1�}���`�n�5��"��@�5;˝�27���YFi�?zn\~e�:0��S�a����y!�����9q=k��m�{GB��(�؀�G�P9P��)����
7�ɀX���`[�WCx!��@Lw�)��@(v��a��s;�a�Ɖ��ICگ<��1�q�6���YC�$lc����d��q����Q�|X,���M/��u5����jt��ރu��j�-?fpH���f���qR���.g*��y ������# �H!��=���[�<L�ǫZ4�_��,�ć�~��������=����/|������b��1W�u��m������Ӽ���"3�\��-��������o���u��-[%�M �& ��R����������!���Ē���yJemL��:&��B������Q��eٙ��/�>�,KQ��].m�x~M¿�#엫:,���'�`C=%�`��MN���5��< ��8Kd�P�>�x���:�� ���F �$RK��S�4�D�I?�C7SD\�n��\�c���=�so��ٹ����#w���t_6���R3螗��&���Mꦃ�׋��i=k�&ڣxG��f��:�,?P���Rʜ*R�y�Y���^Mܩ!�����R��B<�Hh�L �y�mbV�"�B���/���9MD�L����h�y�y����Uj�p�/s�S��G<W�8?�W���zұ}�R�P�N� ����RY�d�m����3lh{ҋ������J��`C��W��f@��2M6�4�$F��Iy#��j�W�je]��6�ǊFr���4�wY���T�ʓ=Ɖ��tˡ�����Ba�z��=�'Q�~> ��`�MB���g,�c����P�䝤qK:�< (\5 T�+\�fE(s��R��`׹��0��BXQ�{%��o�1_K.`/��S�Mf�M�F��\=�]%������{ӯ=��q��"�e2���
}����ܰ�(�*�ʲ�%�n�eDzyV�n�X�7#m�C�Z�5M!�z0l%�����=?+���ֶ�!���ĕ0���!@уwy��`Q�[����
(dKg6qW�^r�2e(ж�8�?���r���Y'��E\1o��=,{�"CQ}���A�n�@�w_�	�e�Z_����C$�G�!h���.�
��V����N拳7 gk\���i�X>G2a7���B�*	���M�� ��_x��/���1��ڵ
��SJ���vu��mH����$��K�	ל��e:%��� Ĭ+d�@���)oʖ=�@zS\��e6)��Q'%h�r:�@���Yo��ڙ�L�̐��/���N��O�X ���_�l�nCu�#<`�ڿ"�Z�N�&��!nx��~�iqC�i���\��[�3��S��˶Cq�:��0Ԓ{��j�wQK #�������݆t�=ɛA�!���;O�����B -��K�)&��������>��e8^6ae�����H}?�,ӭ���?��fV�J�b�q��J�F�W�(���X��K����,�i"%﬐!끨P*���&kG��@Z���u��T���,IP��6�lB���� �@�^G�|�wa��+��k���]�+}��1�(�+e�|o]]���fLa	�"1㣙�RX�������yX��~�Z�#$���7���C��1��t.KT� K�����0w��i�M���8�*@���G�(]�"^dO�fd4�������ږ�o#U�A��&.<�G[�x��U����)�h�� ��d�r�l�2m�̈́�+Y	@���\DI?R��-�d6ٕ�6��!&��m���$��Q�i�ܵ,B��p�M�m�w�F�G���J
�"=d�������EeT.U8q��!�M��0O���x�Dȱ� Bȯ�qk�/��,1�cB�3�C���8(*�z�R?�h岛ɾ�1}�s">�%�e�Tk.�G�.��}������)��P���Os�A��cWRA�����ȣ���t���SB��+q�+��o�g��&�߿w56�%1�Cl�ش$�-Q�n����y�{�`�:B6f5�{Dȗ�<�p4�/�;��`����5ȟ�:"��7R�T���;2j� ���zK/����h��|�(�QL��G�p�(!������*�\��̴��܄��p�ut�r��S웬�j蘛��!�G����I'"�p`�Եaz)���Y�6V�,����[�ߒMZue���]�r��� w���i��=�L��_	�s܌�XLM��	�F�Kp�N:+~F�"Q�O�F1�f�b��ͫ���B���^SB�7l����EC��qw�kOE�pX�N
�Z�w�w!�����>_�)��s�:��q"Io~<������1��}�nNbW;/RF|��|�X�"L�R�G��xϏ�=�n��n�,2�-2L�����F�j-���22u��--.G�>����L� (}���h9��@�V��Z��m��҅�'�u�s̛�K1�<�[�c�A�{氬ZR�}�I��G���O�`�K�~��.2<�(Ҡ�v\�2v�Q'��tV��{w;t�{ؕ��	��p�����H*O����1��:�;��"�x^g��<WD�T��̬%�+9���nzP���ҥM7�=䎣no�4Za3�������޻��!��Dm��"��Y�DX�7c�K���ه�b�y��;2����k�vSO��ĺ�hkĨ�E��O>wћ�/\�"��H}�����3	��6!)��*�2��'���#z=1o5��AU\)L��c["��zP���lO���h/�����H��)�D��*����D��-���#i�Q�K��>�9�V�~��W��\2!@�c��{�#繜�1'n�	 ����<"�A��x�q@~�.i�UF֭���6�3�c��dˬ��˃��-7|l`1���^�B.��#��j�#Z����!��'��eej�r1�U2u�@�C�nM�ɒW�c< �#�{GW�V����20[S����p�q�@I`M~ʻ��H4��'N�0ك���z�;�}�:bt�,=���\�=���0/��0��0����XsV�NV4z5驝���S��YՕr!�;˨��c������5.�CXk?G�Oa���p!�*���~q��,]V�A�?�a��i	��.�&��m�d4��І�Ës���&����H>/6'��>t��&��u�i9<��}����ɔʕLQ0O�]���3�%#�GWJu�"�"���!�Ό�:U�ֲ�'��<4:�Q�[aIj��^=�o�߄K[�G�O�rW�oL���0�h^|�ɟ9N�V��긵f���<�Pv�ùD�.�\$�� ڐ]�q�Ƽ �|�>&bK����s��� W~RpO��{�*���
���o�.�w���$�׀���2ä͛m��D���{|W]�h�͍P���Xg��=��hL�|`X��g�)I��.���&�A;��>١-����(�$���=�7:	���
���խ�e<�g=)�$���[����݉�ѸJ��������Z��Lbb��-&��$��k�雾w@���|�M�B�m�ށ�+;e2�Yu�l�\¤��X��E��z͏H�N�]�!��J���qlұ�����"�Y
W1|:Ig� 1$�&�[�`�ϥj�["��Ӈ���?T�Y�$�K~����`,#܋�hL�%C�  ��`E5T�P(L�`�0��ap�D���h�|�S�k/���>�P��k̝��몰���2.��n;��؄�z��4m[8��$���t�CǇs*��HU���v�P2�a���U��]�'�J#Y|�*��1�I���GQ�⡹�p�`i���=a��f�IvW��'�^rvJV�((�-�\d�������8�������F=�CX�E���¿m�)�ʕ������@�+��gzu2{�m򗅮 ȕ��	�W��^���}��țq-�e��C�~<|��s�=ٌ/%�i��`Z����@t�f+��cd�%1(hI���
��<%k�>�p�ct@b�6�vt��m���ac��v��w�qC���|���37ݣ���wj+�m4|�̆/�[�+[`�m��@bhc [Q�l"�N��w�J9%:U�2��dŚ�����f����������\��eD��r � � i��ʀh^e�T��4�?��}�#[m��j������Bo��M��|��}��E&nx�~z���l%~g�(�� #���� �^:~�|��}��l��.V�[�੡��\A���M�7���(^{10��CU��"�W���8uu,���C�-�p�bx,P��H���|Z��ӥYhӭ�mC-��1p���K	��R�vQ�B��pb���8�;WL�M�BՑ�u��,<] �+��]��s���>��`�U���,�]���#���7�%
%%�H����8�k	���$X�2�#���tQ�W��0Y���xP+��W��_%��z�5�{JT7̂��g�n�ؿ���n�ӿ����onDC�^oƍ�U�(F�,����\�Yt�bt[��d��9���B�<뾕2B�9����ՙ�h@��H	t��O��6������!p�]I\	8ұ�#;�e����~��T7�2P�>���F��E����8��N�͟���cKT�	4]�3o��ֿ��]yMc�_p���Hx���3��;�-2���X�qR:��'@D^fi���?ӕ�7}���w_�0}����v�	��en�o܈��?j"�s.�c��c�2�|�a��ŹK%�F�dedx<N�mQ�U%
�q~)�t}V��z�|p�k���U{*����q�h�u\��|����74)���	�ѸH�]>*q7�b��A}�2n,jW�Sݑ��R�h_6��==t�*y�-���(E����U�1E����ʳJ�]۝�����9��+M�� ��]�u&�a٣�:������bN�B֘�ۅ>О�r����H��W���pn��ަvp�e �E�ݚ��Oؖ�'���l] �̾��Gx��эç!ғd����;�����7$�&=x�Pi���D���)�v)�#��Xxl�`�
g��d�~�����NPl�!���l�U�&m0xq��>�F�������	gƼ�Y-t��itL`訷�0�ףj��0�Yڄ2q���F1LD:m��"�}\�.����*��H煖�
ž��fc�R|	���;�'"�N`;e�P�ki��86Q�#R���1�sZX�_�|]�J�W�� Q*7�1�P��[m�hm�J�]3/�.���hr�7�Y�_�v�s�V��gC�9�ݝ�)\��$L)=�>�Φ��3�DN�Oz.ы"��|?�w��ֵ���Ku,
��ٿ'5�ɽ�_����!�sm\ܰՍ�a�n>�t�c�b�*�0��M����%�*�d��v0�h�!�X��͏W��R�t���"sn��y�	[xs|�2$�젆�oN�@H��L��9�Q�����o����0WGR�2�&��ܽZ$f�A�)��i��Wq)���#�O�@��CLh�_���呺�΁HJSG���n�zke��1��!:=,�i������
��ɳ�)���䪏��s�"ksY,��ꅞ�?<��q[j{톬�|�"\9.M�nZ}PꡙY2{���X��h��l��!�v�L�d�뎚�ӆ=�9��D�މ���A�d��5R4W��F�f���@�a��+|��(+·��<k� I�[~��ʆ��jP{ٳ�+s%O:r˚����%���(�M�����ߣ���>�K�gW�W����`b��ypȥ�<����Qy"C�oH�/�6�������u�)\-;3����w2vف ��xH�ӗ��=�3C��z�'�/��O�����	��.�d0N���}��[j�n���G?����UE>�?W 稕󺁌��o��l`1�ɘ�.�ݍ�/o�;�LѰ���
I%�g(�B�v�s>W�xǇ��8�z�x7���"M�|ķe�x�A`��?��u���!���1�r՝��b���f�m�0z���}@��o�y���~es�#˂}ܔg~ѿ���x�X8��W�m��pՀU�Rp ���L˞~,�.ksr6��Y*��#��U�z���%?!��1��M��6>���\䗓�q��0�G;~����ml���'�_9�����~<]RݸL�Z�j��D��E�
ޖ렝�A4D-�]�j���X�l���7�+���-�NC���	>�a�t~�{P��g4�N?%^��T��)T�F�'2��:�� gF:�����>6��V=�d�X'��㭲3-@9�!ET+Q�o�4��\;���\#4u��?G���Z����G�p�q�|���#��,�Q����՝���A�jvsxFe��B'�a�P 9������U^]�U�.<�P�4�Q�ң��Li�8���҇� �Θ��è(�Rk!���⣄z�;����nU9Ն{���`�"�S8�����F|��͌��Y=�"�1e�H,ˊ������z����lO|���I���߆�s>y���1��PJ�,���j(�_��v�'�⧠6մ5�%xh��G��I�2=�x"Yg��.����5��q-u5��$�|��;��|�տ5��<����8���UHLbS2��A+(}��4����g��ߙC���'�jϲ�l�3��B~� ��\�3��a��@�I�Xp"����U��o�Ɖ�YT��-|n��2�j�}�V�G�S������(;�n ���x{� Dm%��<��}T^�<��%�BG��bVz}��9d[rM`���;y\_iuUШ����a#�u�a��jԙ�����b{�D^o�^C��E�	__�(@y
5�����!���%Z����&ѻ��wSJ��|.�C7�Z��;)�J8sZ.l�s�$!t!���Q n�S��I�5�8�g�^q@��%��;&Г|A��E�#��9M��	�_���T�ŵ�,���������M�e���B�(&Po݀H��~|'հ. u�i%��u�!�6��S�s���*b1UN\��
�s\b�>���҅"A�V$H���i��O/'�	�F~n�Q��+�Ť���z��H&[� ؍԰Y9:��}`��ѝ�pP:�Pmsf�R�}ۇ� �����g�2��^�Rb��!����VG�W����&y,��Q>������r5�*K�f��QA�����F/�!/~J�CPVP�xկW�4T%��{�T�r�v�����?3��x5�z����ߵ8�6�Rٱ$}���: ܭ7\���
�9+�"l:7�N��i���NǅFN��� �:%;$� ,Ti�)b����`��v�#`g��h��eBؓ�%L�����%�] �]X�V;���!�����a*���_|�<Ǔ��u���s�qg�w��914r�I��o�O5q��;-��l������5^��3mI�~n�z)r�0�<�	�[�a�Sv��Kh�9�q����-H�5f��%�A�*�c�bP�_ZX�S� ���B���R?���}��;�'b�ԉɫ]*��b����3��$���QC�Γ1�Ҟ�L���b�kT���	�޽Z7gqT�|�>�j�eP2��tj�eT��=�M�'�5�R�[S������W]ׯ�:�ƅC�B�/���ޓR[#o���ʉm|��4��K��(�VB��˓n�	����pD���J��8��2BQ1���ʇ/#{�LK��Ǔ�B~�O�����A��V�{�	~��X�L���ڭ��ț�%҄A��^�)�����Ŝ	e0��O���p%z�؄�J�*ך�zNb�ԧ�j�П۬�Y��y�.��}�s�n����V�j�ں_i��Js����(.�A��Ve0B��\�vPحא1j=/��t��g��q�ϓ�C�� �'����y  �^�ժ�w��d(�[,�``1�dŀr���A\*0�s�KqnF���N���	��V� �
���JA�zJ��V�`?6|T�@�8���aW���*��{��PUS]���dh��u�훫y�ꌑ��j�Q�{�dy����,ȧ�v�$����$�Q�)Ã�	C�Qb<�{����ˁ;s�~b)���p���^ke�x�\n�0�V�������t7���X\l+���Z�j���(�������<�r��(�)}�cjړ	��5�P"Ƶ2�hc��9C's ^Z��\Ey§p�m^H�bJF��l��d+«����k�xA�a]_uz�Xr�@����rČ��ɋ������S^�f}w�dj�猲|�j��F��x�.��t�Ɍ�׹)$��NP�"���'�;>�ꗄ�1����(��-��h���/���d\p���*�
��J�P�uY~��1�a$���?���ygsl�oa��U���ӓ�7H���L�Q$���5�]X!>� X�s�������DR�dc����~۪�)�,�_�T�0~����6Yv��w�N��	\�(E;ڊ Y:JV%�A��n���vU�V	��=��Z�&���}�qk��v\h�B��Iu6�� ځ%��c�'s�.�
�Yxqܗ�(���)�}�¯E`��H/�O�
X�"V���a��l�p~z}5,3'a� k"� a���ɺ��z�D(�<��8��g�D��|�A���E-���F~*�7�����~�\�C�H�k!T����!�-�r���1����s 1a8�c��';�t��,��@��n�|�-ηB�7\��%�]#&A/]q��l�e��L��1���<�a$�Akqz�DO���^ܶ�����0L��}�g�Ί�Y񽂑ߔJsRz"?nCoLk��wG _�$F��-�_���Ѣ�������-�iB2PN�����9D�E��A���Ng�é
���P�BP��(��������	��r��<n���
�C�T	_�#F��n��QG
�kʍ:/���r�#��D�s-:M� �"���ZFtTN�lH�m��(�7㗳5�[J�I����KZ�L
P�����㬌�g��tO�_I�rZ���v$3�9JAa���v����S[�d��h]욑Z�9	NS�1��)DǗrсz��\�Z��cJ�"Q�8Lw�;�a���N�_MCl��H�,h�k��.��Ͷҟ<���*���<]�o��Hh�C$����"^9�ѰX��l�t��Ac����`�����f�jy��^���|���H���D4��kk����$��4+]��1-־����'�ܤl�!*��K�o�-�J٬'{x}��5����=O�$>i�w���)q`Z��Qwl��.-�O��i/G�^W�˰K�0�0�|o�~f�it�.9c(+�ҭ��u�o\�U�Ч�:)8���i�
S�|��ϖ�oP�7*TSuG���5I^� �c� �{��Zh���T��X5H��[NJD�]
����I�ꕣ@�l:��"�!�_��.�<�*@�u�Ժ�RA-Y���b
$�7"�*3�	(��E�\��ڬ��@�����[�%��FCh�5��l|�E��f�fzO��헶9K���\_עT�u�!��6�q�m��\�g.j�����th�cݳZdl������}+�����Q���|�_^3E&%
���������v�3D��A�ۇܳ��J W88�J���JV��Q���A�����Dʪ0�b�\��-����W��#�L�Gs9ekH����B�ן�T�:�B��j޺��</ t�{.ԃ|C���
��Ó���Ć� �&����?��pF|b������4��<kc�9�_�����zkQ&��[�Ǆ�
�'����8�Jħt�aE?1���e���:�}K� o;�90���yPl�@ԭ����$��Z�z����W�W�iү0J�;�
�NE`>>E��=�����y~�ä=�~���>`�H�XW�x�Q��`pe�a��M�M��x��D<W8�Df?K��AЌ���8iu���<:긞�Z�v�y�w�����)mC�t��0�w(N�3K���
��Q`~��Y'���?�ܚ/�g3�4�(�;8������䗲���3d�|�fX1ކ�q�{|O�N�㉮k�Μ�B�%:��N<���zƽ�W����ρL��ɀgl>�\����2r�������M��S���?@�q����a��	�iȽd߼�h�.�fw�x8��a+'��������xc���|H���X_3����� ��8FtH0��*�/N1����9c ��8��0����3��3ք��b�����Quɒ�,���7Cb�8Ҙ�4�:>����s�0BŢx9�u��%�8JƘ����q��H�}�`�D�+۸!��!6ӎ]���S��2;�q�'���8]{Z�Cz�6�]^�'� �y��]UI�MlDә��HA��*%O$w~�s&m��2�І�o�y�a��(Z�pF�_�I�M�p�*�H�F�k Ƹ���vBe���,@J칋��,�ku�Ǉ-���n�Tݞ���;z����1�OS ���<��ʆ�N�#f�+t�n,Fpm��b��EV�Ok�'��4ZTy:y!f�S9\m1dE
�򇚨�Xi�oW;Cߗt�~�Q2���Ĝ���~n�)�+��~3�s&�?ڊ�%�_t�,
5K���+A��a#��$2���I�+!�l�I�,���<��e��*�6�����\A'3a��؛��)Ք��tJ���Ѡ:/򛱑nɪ�0��1	��E����'<�+/b�����<��F�6�_�)SS��&�׬�P��w�zO[�~�\($��T�x��5�1�$�\ �c[S�vҚ������[P��Q��=�pNe-��J�x��köEʮ�����q��~�k�d(L���̏D��n��ϵ�v��g]&�IU�b!E�0��M����8L��h��u�J�j�j��eH�����׮kjC�4�XL�$�P�#�,���1��,P$�ݸ���02tt�X����\A\��6��I���H9&��."؜�����yMei�O��	��z�K$eR��t ��g�3�qB��H(ȑO!h����	����Ȇ���|n)� Za#�y�=P=��|ljEBGƐbV26��)�� P(�}^���]5T#��b����	֭���s�� ߳p�G����fI�8��Y~��V���D��I��?�ߋp���M��g��x�a'��Oxj�����v�'W\��#�Z�u
�gZ'�u*\nX�k���̢S����{����!_N;v������}-���}���C#0ov
{H�]�w�u�s �0�d�H�E$JH�]��-H�3j}n����'�;�C\�X,�A0	�5z����� �k�
p���3O�'D{,`�f<d�!�i��U����T� �-&�I�1b���!^}D��)�|�Z���{Fltߙ���i��/vJ�߫���;*�����<>��E��t��%��p�EO�s!��@Ě�*=�ĥ�W�؄f~��mv�!���?��/�/�����S+7U�p!�]z���+t��5kf�)����w�ޤ)�w��t�����?���2]	�A�����
�K�V=
1 b&h�h�Wp
�cM�o_11��'�igk�|9��(��K��0�A�2D6ȝ��1�\�֌H&
qQ !i*���e�WW����丆�7mh�'�]y}N���"\�w�@1ƪ��?e,���\u?�΀BV��(;�RS�n�5�V1(ȧ�GO?�a׺kYN$��C�7��v�~����0�7�7��>M�(��=a�(����m�U\$.`,�u �h��� �d��_�����t��#J���`-q����7绹o>�MYj��-�=GP�s>D4����>1@����խ�{�o$]�E$!��]	��C+&t���I�k�����;�FW������F��'���u��ZMO�).Y�
�F�?�`�'�gV�Z
/�`}�� O�{ށF/��Bs��dR���q��սKl����9�J�Z��y�����"{[ēKT@��z��}���
I<ձ���]�������p�h.��qR��ˣ���~�l!:6�i�����JY�g��U�����2O����s@��"��pa9!�xp�<Gn���Ǟ���m��`��I,rԸE��_����6k`�s$�U�
�G�����T1k���d4:ȃ���ojݖ�4�6��(�x��>GKH����)@,?p��j��=�m53�.5���U�5TQCd82`̞]�&�;�3�^�i9%�+��
�wQ5��s�c��D]�U��)��8�"r�v��`�ل)�ݕ��8k��YO�I���#������<r��O[F�P��J�Ep���`(��+�AX��C7VC���3!/��="d$��r`<�(V�M�<b�cP�gY&�S����z�M)��b+9w�j�_�-���-�!�\���W�����nd�ELEuW�6u�7�6���p^$���H�o>Y��rLb�|W1b�\���'���r"�%����v^%$�D�`���BW�?�ݯ.�,b@u�3i��׬��Ov�B~�t��
1Z�����un�@� �a�/��%���zMͲ��.��`+1R�~�ZjJ�KQmi@�ʫ�}�l5Ϝ���	]����X�$��T�v��vg���[��(��$�$��lZ���$�b�E�C!�ƹ��%a=0�qڭ[�k��S!�u��#���A��q��
��%M���˪�C_�U jd{e���z��X��9v�	V�F2�}_H& V1s*���3-����Y���MUJ��1�J�u�k�/br��3���
�ğq��6$x�kx���J��i!���Y�DVpď�-&�k�{�)�J�W���KƮ؃lx�[�h�"68�=K'=�0#��5o�6ے�I��uq����Y�f*�SNHϗ)ˢn�C	� �����sd �l+-}���Ƌy�S}��]e!A�0��7��[�vS��Dp���Wz��=I)��MD_}B$�<]���bM�{)����m�a=Ğ��heN/������;���� *�/�HC��M@]�؜��6�<58���<Ժlfm�h>�VG�&8��z�h"�s;�h����Ȫ�5TW�_V�������-+Ó��t`W�͎���$���/�ݥ�$�|=�m�k�iJ�8W|[���#���"��$����K�YR�)
�w*6��բȧ�y�������2��rn4+ݶ�����Է�aQ�1�.-�3 ���O�UJץ��(OY�cƝ�o��$��)�U��7!���А���$~�2�ľ68M��f�eR�~,���pٚ�/�H��>�@�G:�CW��PqZE`�}B�	"�qH���fm�,�AAtc�N�'���T�s+qR��ɣ���8�w���Ֆ�3�ّ%N��l�����l�1�g������C��3޽:Qk�Lf���n�y]�J}j���h���Da5u<��jF��EȰlȠ$́ɼ��+L�_)(PH���Q�ڗ��x G���������rH�_4E��Vdr?�0�r�`QI���s�kp(��s'�,�Ǒ�w��v�RM1��?Ȣ@IR�,J��oo�35-�"&�gy�E�H����)��2k��kW��˵M�Vă���o��2��`�/���A����)�����"�재���I<<�vp�T�)�l�ɋ/�Ĝo�y&]�>&���^[Hv�b��8V����{�n�qy
��Sӛ���>W����5�aP��Y�t.G	Rw�^wҭ���1d��v��'���^����=Ov�"�I�6�m"��2C�_1��[!~��V<���h;$�h��I�����X��'�5��x�xe��Z�ωrTǋ0|�� T����_�y3�)P�l���f ���tC�]����6�V��Y�T!"8��������
��B��meKs��kѤ�0�n��ÍpQ�2�M���c��eD��#�H���W���d ƇY�_�����CA#;@S�p5`�Ш%@�W{7MW*}EY$'%+���	݂N��x4��DU��M��E�pk�k ��G$vhNRyr�T���#���TA�`Km��BM��Uǈ��T�~Q�Jhg���&sQ�T�j[_��X���?:�D�+'G��I
�A�0��/���f�v�xds^ց�Ȩ��ɶ<f��v�7̵��A�"��!�U7�z�adR���lS ��ܧ�s��F�ON�*R���5�Otڲ
*Z�I�f7�ڡ�Ĝ��_{�F_|jl�UoRM)�TJ��Vb�W\gL{%gqv�cNSt��O����>@CГ��N�����U��)+�*;'
�V�r�_�Қ���(ۃR�y�4:��3�<{cOG�/6�G�Y�ѹ�:��C*�^�@\�y�7)�����Z������h����1�،��@�D��2hI<���\n8<0o����w��W���zG�k�gp�,6�]�/��$����>��a� ����Z�s�˛3������G#}�A�oGZ���q(�# \
,���ϟxo���6!f���(���Oit�WBxz����s.�ҿ���H(��sy=������.Տt���Kh�
�C�c+�򙶲B�{О��8�9yT�����Jc4��ڭ��)r��@��<���t��#�8$� ��ر#��]�Q����T�k�>�
ʒ�D�~[�r�A^������ay�B�(͍��)�[��ұ(�5�t�T���zX7�ޗ�#:����y��"-�A���DW�4�΍�o��Ҝ�`8�U�P7�6���U����YK�4�Y� v�����6�!:U�w�<��K�B�G$��S����⛅�\�}���l&� ��"M5����
���Mq�:�b}�K�	��Y:���1������\ɶ��=���h�3��ӗb�g�a�@y�~~�Q�3�js��a�QBX��U����0��X�i�� �.�y_w4;(���[��+�t�-��>Yg{�V�T[��;[�eꩾ�|�>���&<Q���#��?�\�}b�v �8~W��!�7Nm|ā�Up�%7��U�h��)Rx�!X<�^��ըi4�og��u;�]ֈe�Xv��Q5�cYG�d��"�ކ��D��S{��GOo߸���f�p��[pk���P�h�����&�G�
Qxo5��M���Y:������h��c�
_��Hnc�F�ř1�Dɶd�Ȥe�T\�|��SF���؅����
��{e��g���fb��;!a�d*��פl3���: ���)Y�t!����c0ŴQ>"�jv�F3����{/��sMЮ�!��������ş|��������}�6.�3�y��52`�m�\��
bj���z�I�� $�GCq�A���k��:8%���'j�e9�AW���`_�uվ͹�O�o���>���:��������0dB$�.���i�Gt%�U�`���WL%��X����n��)ѦsOf�8��Y2��(������z���(õ�*��y9.?_�<J�� D�W��)ݑ8�
��#�e���k�Nܶ@�N�'�4zHy��G�8gRq�s���Y$ �օ���yڧ�v6���V�����0��\;�]1���}8.����P�@�V�����-���E���yf��5����@�`��0=�D�"�0y�4P-�9�`�^��w�v:��9:�,�|xd$�J��IL�U�g��DXP�P�th�B���J��u�V�Z^:y���B�� ���itos�吥^��d�rLą윱)���%R�)��9R�f���6[fv�P��y�F��;�Q���>��
d�y�' %�P�Lc|`ӼU�s&s��0?9��G�X�"r��,B�Lp���[�o��A��1��m�&*��Z�][� C����U����@a<��_*%�c�(zCǯ&*~��2I؏���َ3 �����:�Y;�:�;N#��n��`W��䌦�Wn0E^�����20�����&�#c�B��p�@V8�t��qq��� ,�T��x=ֆM���nɠU6�\S��o�R�'��dA�G4�%Y�8�Cן�͸�� �T�־�0V�NE�Z�˝ĉ�!θ89e.����$�����L������@k=��z?�ػ���}�� 
�-�F+RmQ1��́�	�A�X8I�!؇�,aJ}h#����N���?��󭑓i��eز��>#�=�f���n.�T�I���3���o6�-&���L�9ޤ���j��ie�� DR�v`����rҧ�����ج~ ٸ���$��Ž�%ބn��	P�.Ty�=��S�~��0��:]�J�f0���1���etZ���I_.Hx(��ǥ�,Y����O���K���$I��ۭ=_�[��AUܞ�}�P��b�������/8#Y,�P-�0Y��Ѐ�)��eo��#wg/����"�u�O�Y�q��MXЛQ�Y��1t�V�Z
�׃���!�J}��@}��		�ヨ�ʞc�n��-�Fo+�w9s�%�0	�j�م���]{D߷�J�戓x�	��R �P�ߢ��ˊ����&���m�-�{q}Y�o�*�9�Ъ!�h�3B3p�uN0Y�
������g��f�|�O=Qsl������*l}xݻ���,��`�R�,�,XQ����@�ux<�ܱ~���T�7�P��F����-"��9��*Xe�/�R�t��_]S�5aLx7��>�v��]�ܴ���@w�WR��óZ4'�	f+j0o�*n2_r���D��ǁ@��~��8�k�ul{BgR�4N�0�=��s�h~�WG�p_,�N��95��O|c&9��ڼ�0L�ĥU�P�WԻ��\�����������a�{��6��z��o��=�$���*1�j�=:_i��Vj��W�,�l�!{�$+;]�2�ZǼ�p^�&�չe�q�PIh���1�[$�-����h40y��>�Y;��5�XUN�Z�sJџ�#��#1��������9g�����K|�t�_b��ؚ��z��0-4/jx;[)��5��jDc���^Ҿx1�nx%�v�p���"?�v���zߟ��*Rk˚B[��FBU��Ͳ#S�RɊf�Iլ�Z=@#���mD#�ҴJ�A�
���lM�of:!؂�Nx��u�]�ǎ�](f�_�d�뭈���%�8��O=�<#�Yd�D
-3&����#K�]�x��p�y�a[,A5��`Ɉ.�M�ߜe0�mʑ[�ʗK���g_�׌Z����`]xm�����N����{^�qH��'�b�B4�8[��L�����Jw	栬��o+�ؠ�������^ù���2ư��X�*�T$�b�W\/;�$E�b�G�~9	\���
�. ��c���`c&<{p�����*!�Tec���'4����9|����>�!��C�(�ҭ�6
9����r��V@��b�ʊ6��AoC�^a �v�:[ ��F��x7��0��W��SUP{LTN��G6UQ�b�����F��7#lYֲ5�WL�
�������]���q��?U&?_a-rxN˳"����`O�^���i^"��ΠW�v�#�KNVP��.*�� Q�uc��@�V�J��xHyU�뚹��B����+]sVca]C�&�X���Vhp�y2+C��B&��m����;�ld\��?R-q��ӣ<�U ��d����%��<.%.����7.E�0�0Z�}�n,�P�������Ϣ�1FctMj�i_!�.��8g|1?Lm�xf�9r*����97�2��/BΊIO;t�&�x����T��҄w�ZC��]����D���h4�-<'u����t��s���|���s�,߈�"�Q�@X��g�6�z�����&HLW~E���,�:{�^w$�
��{o$t9��C"��^ ���!��3l$��\h�
����3�c�b@�����<%
>:Q75;"K�M6�ː�w{h�����hD~q1��Ϯ�3e���E����}�g���!��e�L'���d��y+*+�s�^�S���n
��i��B��ҡ�<V���c����oud���z�Y$��>G'%�?B�~��N�� �q�7jh�VáƊ�A)u⋳L���m|���1����s,�;�s������S��2pL�M�q��s?����Zj�D��Gf�P]#o�o���Z�����:�(���i����W1��%<���3��<�:b�9f�Ci��ڃ�A_��(u�C�8¹�B��J�QJ��'I�E)2�a�O6qj���=��b�9��,�Y�6�9]���T#��>�n�����SA�)���be�A�}�H�E`�����&���:��9�ߔW��O���1W��d���K�����l��s��/�[)�ޘ�߰�^���f�O7<c��7r�K}e��{�p����G��!����ç斜ת���.��G�3�pS�>Q��(#��h�ESRͼS��V ܎l�N��V��;���nYJb�_�%���6�=g輀��&�
mDB?��]��&	������/5{�./�q8�-��\�,�s����7�A^i�_��bN>�p��`��7�Z��I1�X�9Y�`������NV'��?���J�t� .�Q��
qnt�z��8GD�)�/w%Ϧ������m�O�N��8�S-D���(�SFQ	B@nL�x�`
��g��B}�j�^3���"�F.#��܍l�K�;���x�3���RцL]�n��8�E�Vp*�=�K��u)D�y'���h�s�rXF����3����W�(������e�O�� ��OQӹ��@�e�ϐ.Ou��K���J�R��C���LV4�6�MД�sP���d�Cq3��kc�g�B�&j!��5���A���I� �����[��t'�f��)�Y��a^���>�s/�ǈ�h(`y|�5�U��Q)/U���\Ym��>�
�G��@m�hq�0�F�s	 �s�J�u�����gp1,���4N�ROl��=���۲=:����n�'5�������J3�BT
�=��E%��:�����a�QK���Q�C�8�8?�5��h�����w'�K4J��+�T����1���#0'aV�Sx�dE7飹8�Q�dS>!���3���^Y��Cf���ۍl�S���,��L�Z�v��4=0����!��m��1<Ժufg���zu���?_E�V3�|�WJܫy�G�GE4��	��b�ˈ>�[ȟmK�}�Q'mo�_Y�>�aTȥ��}�)͉���KR9�tp�8<;,��tp�w#�S���"�|z�(�Dt%�P9�[\�dbBI{�-�rޛ�����^E&C�H��_zk?�{j�퀑|�qA"%���q!�g��; *���:yπ��5)�/�|�^A6��DN���r��5.7"W���@���vg�]f}Vp	�~������MH����V�v�P�|�@��z�]�+[��x׬��#_��:��Z��.��.�l:r�rx��y}�X�ŵ����8ٿO�0����0łsx�'�":�YJB$lmأ��9?L�y/��I;�l�N1�~���h螆X��كOW6%4����# ����k�ת�A�X[i�$��m�a*����;w��u"��W@iZq`q-��:�O�ށ!�>�N\Q�����z�8��B8��k�dg�k�K������#���JI΃����	�X�ߘ�e@q�	�� ��wg��� 䏮}k������F�79�]�-k��DW�hS�	�q��/�V��/B9^V>'@mb�D���y�S��q���x�Ԓ��.����ك�ы�X�I�q6��48Q6jF�Xߟ���w��,���"\UN$���ݱ��|���d�2�m�+7�O/��Z��}0&�!���;$6e����`3�dr8F|H�W��yA~�W��(��Z<�� �����	%��������~����n�mFGZ�fQ턆�w�?����c뚲��L�O�^�~8���s��s�(؃�R@R�����S}^ǰ��z�=HB,4�"泟��uv2�@<C��(�����[�Ppo��0��#�>�����,��z�S⎻�B7�9e�S;�qV?1l�hU��7!:Q����Ҧ�o�C
�k�7U6�̟���W�9����i�?hb��l4��q���"�׿�725������]L���mLf���c]<��P������[�Ű���m��D/���>��}��oUB�G�d�,�QY}�uo����\Q��<����E�N��Sdy��Z�����f \�,5����0�B�LI�n�y'y�	%�B�,ޕ��{�|z��O�0���`*
W�؂K����M �������-m��ʰ�j�S��� S����[*������FT��/�ފ�0g����QC9[���"
i��7B�K��6���'�<_�كĨ�A	���v�LR5:�'�i��.�0-�:�\Q],�R.ư�hU����-�ךĽS��Q�J�" ���l��%xا�[�.���Ls�������8I~��������A�7���A�К'"�|������l�T�P��\���%�Z߾�1��HZ���y�T���|Ռt�ʼ�ӕ��(��0C�B t����jP�2L��}�U���J��I���:
?R\��Z�`q��(�C.Ajp���XBr2��`J�?�Q]�U]@>���;�.y=��_]��a ��%�ua��jm͟}�3z��iR��]�#�FE��)m��	A't]V6ؖ��t��(V�P�:��{����@Nk��C�k��.ud�>��Wh�mno��� �OKND7y���L�D_��b��8�U��r+���A�϶���,Ec��k�H�P_�]R���{z�?n��j�@��È3}�C<eT�	u�G"�Z���|*#�;��.�V��8�4\�v���-3�S�c�Sl�U�"��諲?��0`�\U�bV9!ۅ�=�&�����ŀ�ϧ1�;{���y�J�1�j{(���җd2$[���99xNa�L*�v��}���d�+ �y�E��+����08I8Ekr��Ll��y�ro�? G��zkj0�|�L��a��7�lnX%/[��3Bs������S����|�r����M�7���֨���؄�2����}K��!�e�f��#(@��e�fv���ϕ���BqE�8TQ����,=�I����x ���t �9&����+Z�J��)�10���p�C��3�c&��	�NqA��i�R�A,�k�10C22�m�],���
D�)_=t�k2��w,F���C�Jw1i�Y�_�8�	���R��E�[�|�ceM2����;��2!-oXu"�y�aչ��D��:M��&h.�6�ӥ�%�*i �Q}~Qu��PR�����kXO�G�4��*2���!?��q�8�3�I�=�z<���qP���i9����/��!ؘ8f�#!J�����atx���%�4/UC����1��2���e���1R>s��0���x�Cm5����4ۨ��u���d�Wօ��@D`-7cb��*�#�3.Z2�^���Sр��)<���E�夑��l����;�����Fs6 �ĕ��Vq���1F�LS�w>��o�:Q���ʆ�%����ʈ�j��W#�YLH ��jD�-%�ֺ�H{��r(�e�5;�;�N�Лp1�ec_��9�M��2SϥֹM{���MTI9ʃ����dS���T�mlǑ���tk@��|�ǣS6�ƥ����dƣ�#|k��on��I\���&��-`2�1�������s�t�QSuz����vXK�c9�6*�UT�K:��%#2�(0���+�o��]�#I�P����"�R�h.+<3Ŕ5�EC=Μ��TZ\i�� u<�p�`~�g^e�� tRX�l�s��O�<��� ����8��Wy u���(���`�ׄ�u�+s�|/LNv��MlB����B��'#]��.P����Cy�8M�9�����NxV���� I���T^������93~(�8<�="�r�JV�z��}�;g�E�-�1f��׫CK�Y�D��[�G�` 5�	�k�>�Vcl��s��(��k����J�Rͫ�I�D�ߤD�:H�S�� ��`�}���j7�n��}
�p��j,a�A�
˲T��$����+!Q?L��[������x��,'�9��G��9�,�|c��y�+aX��O,��������\4��+�w���XI���Gm!�!���
�����Lz��^�/���0=oQ	�;���'GU���'Z�5�B m��Ki3	���H2��p�+Ʈ�!�ߘ���*��S�O(���q�O�s��+F�'�. � ��g�q�*� ߭L�!j�r�^�:�G��F:�0�����V@p�3�H��9ymY�E�GbDZ��)�Ц���e��jA
��)��ɍR״N�o}����[qf�/�/�ăW�[W�2]�\~�/�J�w�c����N W���̼�;��F ���
=Tv�<S�&�CY�a�bNý%� �r%��������!��� �)Jb�;h䝉?��a�T�jj�13����i���U�x>}�/��؉(�}�@��p�������|D~�vGS����Z��0�W�ft,��z�p��+U&��?f1N��\�M�(�W����
h���]4v㷴FӖ
��H�0���5��#e}@�h��4��v�Q���J��V1��}R�]��kc;c��:a��3�X����0Js���sz��fX�%�B���~5C�v�A�*����F;aA\���yЈI�g}��tsZmu��A&��R�D��F��ĳ�c]'�3��K�	#9v�t�9ˠǒXŖ��g_xtǃ��7}?�l��F}hjҌ����e��FR��8�G��J�Z���8x|��__6
�~�:J������`6⛩��`2k�^�q@�`�3G���fp���r�|�i��������V۵Nrb�
?-�CG���>7���������De�/�J@� ���ԅ8�D��xsW�?�Bs|���X���|~Y��Hx�6�>Z��g2^b�����g��\�zje�E�6_ >��L�y��
_���٣_B�r�[����1&��4ZS�0AɫvT&��d@��GY.�'�����	��Q��F�0|*�$dϟ��X]�Y�)�?���VgVa�`pL�WL
�`"���6|�R�13�F��#�U'�R�b��i�Է�S��yy�������A��n�6RJF�4A��(�w�9�XL=Q��Ƚb��|-6_�x �Ȭ_��Y�B���_�,�0r��ê1�N��u#
v�<Kg8����׻��=�����ʨ������#��엌٫�-3���s��]��;w�oRy��Y��������z).U���e��ՠ���.5�G��5L�	D�ǚ�)�ԝW�F���):� fE��R�R��v!/O��AG~c@ʹ�ן=�Ȓ���*��ͤv?���$�|n2w�P�ky7�yF�|���G�(g�C�0
�Bu���Ǝ�����7I�+�׌?���J&򕷣%����]�Bd�<J�ߣj��(9�h�<Σ�k�m��]-qB��F'0 @��7)����p\oqI�����kD��֒��/Bo�{�Ҧ�ʉ��@��QD�'��cA�U.�r�M�qFdS���4c�*�!v}e3�'C��wi��ȁ�Kb��Y��T�W�^t����#]IQ=������@?���V�/�.���2'!=%��2�g?43e$��6�l.���VO&ȉ��?W'/�ɪؑ��ox��:�_�l��G*a9jc���Cq�Q�{��vLT�F:�1z��}�z�kO0�d�~!��r����ǧ닌�D��.���7�De;��e��{��c�����l���-��rQ9�(�Բ�t��g���%����A>vF�����*��5�؀cf��.��)&|<_jNШ�w����lW�nr�ئ{������؍���(޾]�Jd�"�{L±A�K|�����"�!-��Q֋�-\	꠯W�����9�qJ�c�3"���~T���m����K��4[;���l�G��(���:���B�&w�Q��{��O�a� z�?|\�
Va
0�+�'�ܴ�"W8<��B���̣#��t�=(�T̟���`̶�ɃN>��׆R rI�dߧ��&����UB�y��=��|u��Lw�ta\AC��8�����п��r��cLi����8$�M'���6���!j�S�಼>K�YH6+&�;�"�P[��U��,�>�!Q:�0�=E2�����4Sd|$/��>o���(6�,kh���K,��%�I�!ZQ�	�:��BN����� >z��j�#	��#�( `��#�-�8����gm��B��ZT���`�[Չܹ+O��X�Y�F�༄�
�}M�z�(<y��)�&��_����O-M�e��*�A�ߕ��zmwB=�m�W�B!]9�|����),򺓷�.�ؾ\�\�^��2�%�eE��`=g��J�Hw��'<�_���D�Q�h�<&S��i�fY�����wUs,��8��[��|: �Ԡ�$�v����u��M�Loѕ��Ps���#����b�IL�+�ƽ	k��N�ݠ��L������ֶB-��x@M�{%�T��%�������,"c��J�Kꨕe���N�3A�F�,�2���|UX��ɬ��~KSrc��`N���X0��Kp��J������*7,?���+-�>�b�1bL�+`�������tyB�����u	�홧���D���g+��i�g����10�!�R�����n��~zP�S�А"2޶�n�7F�z��ʠ�(��x.���B�򲱄���6�)N\�Z 2�_����w�E�濚���#��m����/@k��C��<�w�>��H)Ƌ3�hc�l�s����4���n�������!��X�T��ym��H���J`� �^&���)~�ZN�&�\!t�O������e�S&�8��u,?���O�)N�D�셸9E�Cd�+'B k���t|�;p��U��5��ߜ��ɲ���S�O�X�0�khD��)�������;�@ZDj��<��Ĝ/��!)e\S+�7�35#��XB&���4��T�H��3�?��o��>��"�B�����?4�I��p�%(��F�ɾ�a�dm1��?"Ǜ�̽L'�ݵ��a�^�u>�W�N>^�#�Vc�Q.p1_YȲp����O���U��f��>��ٯ���i���;^�. #g���'�"��fjdH���<�b��.K
�QZd�W�CZ4<�
�ϡl�ګnD�igoc:�*���o�"��v������-(Sp����/��
�0�^��c�j���B��9�ԁtc����oEYv����jP�vM�/<�ߊb������G}%��n��p�]Ĉ�����	��+KUk�s�� e���2��<��eE�sw�J\H�ο�2橪v����c���x�Y�ύ��-�ݮG��d��E����1���Mڒ�Y�Xa��]����^����X"-u�>��$�#��]3&�!o�A@�j7H,���س�(Y� ۡ���_Ē�WX%�E�6:�R6&�	Z��j5��g/Y�vp��S%˕�E�z��,�C�a��1*;�$l�����aZD=��JA�y� W��c��?LNi`HjY����b+W�i���6(c"�.�]^/ӦͶX�����\O��bw�L�XA�����S��4@{�w��g�p�y���E\`�ΊUؕգ{8L�1l����!�x��A���*���O�_ǜWGKqj��q��n�j��]Xm�7A�$B���q���v�qCK�t���s�)}݇��-;ñI���+vY�i�ɪ&��
�u`��|��g�l?�a�kK�e��J�������/��kY��43I\C���n�er����@���B-�e��^�(-�B�5]�ژ��"%mzSv�7�	R����q��&؀Y �����j����)�6%�a͢����{�ē�e2­�J��{�Lڔ/VZ�q�n�ˇNx��ݦ��	�N*�r8��\Ar��ء�b����m��2� p�H�Ys_}̽:o�N$�&M�[;�@[M���c-�k[�1ꓴ��!5X
���ѹ껋���{���|�@��cJ�a��Vkݱ��<b���*/��hʄ䋾_W�f����fg����H4�ڵ%��0��I2( M�\)[$��� ��D���0�1�(]�b�k�2�^�\��o���!\ҵ��w�z��Һ��x/������}�Ye�wp���$]�o"f��VH�M_.��M�b0֦�&�,10@�=����R}
b�Y�-����0��|��nB;�JmR���+�!���45�F�� �������'��=�����G�8W1��ҭJ����빆�`R��R�kXP�a�/��k�>���D��f�R��2�K-�O�S$p����72��Y��a1�d*BC.��PV�����@@uF��"��⦏y�Ɍ��N���U��D.%����f J��t������}Hղԥ�.*U)��%_sNe	69�0Otܓ�}��R��o�_� �W�c��KBD�N�I������V�\��(ک�zX���j�g���P�
7 �(iҿ��3��l��-X��ê�@.�} �Um}��?%u��o2�l��#��-��t�Γ�%Đ6u�>RpNJ�	Ö��z��ic�e.��n��r�ƌUC�D�nUPzl'���2�ݹi�齍Fݮ��M���8O �c�:��X�{ �t�[�9�Ag,�)��A�H��X,������;�7~I2bM��Ld:]�qe6�$o�2����r�P��U|x����+����w� �N[gL����#�R��^�?<��s��#���5�c4q$,�z uI
�o��� n�#�3M��7�01���a�02A��)�c����Ԯ��Q������u�L>!ۭ×�9��m[&�XF.�g$^6o1�M���v&0��)D*H��B;Od 9�5�`�^ �d|n� r��g�"{� �m�v
Dx�UG������/��s/�E� ��]���u�rE@q�.Y��p�~�0�֫ V=�9%�v����
��yV�.1�Mw/�@�M���!t�����^%��O������;ӫǰ�9�௻�|�0P���nV<)�����B��LPL� H�5�\��k0�<
J ��JH�w@��Ww8]���2��񉺷c�[-�E=�Q���s�ͣ������ߵ[x�Sy�hΞUC���yA&֟��B���>]��I��XJ���\��!I�D���r2�@7�_��0�#`W��kl(�])y?���@�����7p�t�
]�W���t���{QVα�Y��P�~_�z٭�e�nbQR�����Θ,_���V*����<��- �P�?��7����f�TAoK��ţ'��u5� Ef�4>�v�\�~7��#{��q�)�d����F�b1�-JYri���V9���C��f�b'L�~�پ�B*�u/nH���;G����G\~�;�$��@E�W�83Q@W�H��<��Y�J�a�K��;�O���4z���s�)�x�~Ŵ3���
��?`v��2ݘ�VbϚWEӇ@�SX9��I���+�Ƥ�=��p��z�qIa�ui��i�ۯnlx���RXi��M�8�8�LU�����Ç��nͿ�CYM�7faG�Ns���$<�mtwD0�i;��t���I�9��B��4S� F��[��'z���-�|
�ڋz?+���!Q�P��9���~N/gBw� �p�L/h�^/y�U�9i���y�c��&1Β�YD�
�̓��wQ�_s�0CXޓ,�̪��j��`����>{�z�݀ؽ������c�݆э�����k3���E
8x:D��iD�Ff���*��S���*���dx���Fb��F�VWP]LE	�k 
��b3�����x��e���F��RF�n��1Vǣ 2[��J4�Ռ�Ǩ8 �%m���M��:V��A-��ʠ�}�� ��\Z�ઑ��<Q�g�8.[V�/�I�rMT@аys"�b����@[G�¬�v��Vlu:v�ز����R��	3* ڲ��{$/� ���(�!�|�BuZWk�!���b�e��H���Ǘ5h�z��dA��ܻ��w�ʡ�`��Jê�g#����q��Ho�PJ��f�E"��j4g����]_;�Ќ�yY"�S/�K��Wn�l����kh�I���r�w\S�Dd��-J;?�'`���@ܺ?3�×����u�Qk�1��U�fY�m�CO�_��ٖ;�iB�Ν���ޯ_��\Gd�4�}�m������ˇ)�+	\(�ܠ��*pbm�����<�LGɓc�}���6��'SD�iD� ;)a�_��jSzG�X���aO����$fAF�l��&U-{=u����\Hտ7o��h>{2�3��	�f�������_*npC���w���D�?`3K���ۍ��5�B�V-_i�aa�_���2og�L��aK�N�l��V�g_���=�Lաd�C��8�:V�1�3S>%��90VV�zW� ��=���~���
�vG?~�&>~����GǯP;����;�B��!��3���πp�v�P��^�VωƏp��%�]u]���~ء�(��a]'Č�v���\�%F	+b��d��?7�e�E�v$Ο���kG����O�O��� &h����?/������:�?/���Y78�-Ԣ4�-;����]ȓV)�ct�Bo*H_K	v�P�㹍�pF��4�D���[��i/(oݸj�����1
� =m�����73F���Q'x�Z̫r��D�)�����c- ��#I��M��Ø���gX/2g�y�����{~�����YT�bvĲ:����V��ח&9V�i�z�'���� С�I��K@��ty�Vk���)9Ǖ\C�e!i)�+��^~�o^ê�d�/�n�0(�򩽥���V��f��pv
ȑᰇ�u�D06�ط^8�ޙ��>��(�?3�H�zX�B���t�D�!�ͦc[_h�'	Փ+��*V��ϡ��b��<�8�y%��/��"z6��BF���Gh��D>ho	���`��wj?%���Q�P��Df�8�����Fbɕ�1:���=gp2�Ӷ���l���U��uk�,���4�QzB|`{��`'�'qt��ޜ�4��9��(5g�ȏ�t�ȴ��/��m�Ks�������l<+" ��K����Vm�a��&�}����x>����E�"Sw��KVԲ�M�/lv^�|+y�=��^� �]mN�wi�q��Ϳa�i�HѼ2+�e��c�YIj<�[�s$��K�1uӠ���
_Yo2���H�}��#u���a���}{)��l�?h7�|�D�?<[�I�D-8�M�00-�ם�
N����*�%|�_� t𔘵��W�D�!{76y�2���\��`��gB$��Ƿi,�y�1Kd��~��3a�k�3Ĵ�t?�����C���Z)ځ;�>���Ssͤ\wsd�PR�/L{r�I���_\�2��)E�M��E�)g���}a�9�W��l:�eZ{F��"�A5�rA� ��֞q5�J\��HX���e���O@ �YR'\��T�6����N�[���;��*�Ў�s�N��4���O��K�$uW��@�e���o~�䌡~�U��ē-�C]B#�F��'���Tu�Ucƌ�i�F�Q�85x�6�^*
.�o�Q[������nN��027� 
��a�F��u���h�&��ũޏ�HE�?��m�����Q���h|q�|��(*�h\�u<9v�
�RE��F���ްZEؗnXΘ�/�\��A��G�y���9��$�ݚ�mva���Vk0���s�x"���n;��đ��,���5o����]������"�VS�k���Y.=G��=��������3�������x�Y��9�)o�O2��Tm؅�.��q�	���և8⍲�y}�D���9�S��hp��vo��mz�7��W,_2��!��cR~|q��w�^�r/R�Vu�\:�Mn�z����0)?���~M���_�'tb�oU�y� ���+M)p�/iav�.�1� [\�q�����5���榫�t��Kt
���V9 }[�W���0��÷GlV�����K�̆�2�^�ln�TD|��cqLr��M������`�hs���Ԗ칦���l��ٗ�����m�"����1Z�r�{�b��Np��b��S
{�Y'�PK���?�-���{�.p�� P��aɲ�&�q�)�Vt�Q�!i 5'��{���˃'� �.ݏ����N��m����z�C�������<:�[&�>��d��S�Tl��x�@�������*K?���f �`!S-8���_�Nޚi�д�����O1��Z�U`��񌱈	��Sȫ�da0���l�G���4�r!WFH�Wސ�!iޓ.Nj-Yt��o}� ��Zy�+�Lp�'i.�6'����Ξ���I�H�R������S� ����A��dz�ȇK���JF�X�O��x����۬Zl�{j��b�m�}��^�ꜧ_�mw�I�d�8r�����muV�'5�e%��z"�d��w��$U5j����tǑ�������/�V4�PN�+ƚ��׫i�5��L6gm<�X�������_a�����#]�����^BV����G��(����`�!���.S�����;P�DK�9�U��8ܯ8��
�J�\�Շ�d=�z扯Gd]�ġG�/��Q04-E䷭i��[�@��8� ̱2��O,�e�g@�q���`ⳣ�C��J��A�Kg6����M�JE���ׯ�Na0�r��]��ߑ�����)��,L'J����6�o�U���v�,� � ��l :��y0(<J�E��[��v6M��W��oG�*����0[׾8C�y
�����:����t��5�N���஡Hp`ج�Tj�o��i�����3-|�ײ����H�w� ǾXz��3�6���5�F�P�}�d4|-�;������&� ��<mj[�DT�$ܾq�uPco��5�m�ie�XU΀s�պ�˅���@�)�)Zsc�+�me~�^:K���p�T�p!�}Z��^�1�Ed��5QwX�m�f��������~��d��,#)Cib��4/䟵�(#Q����hr�
o��X%��|%�y�Ǵ��]�5�Le'l6��T�AE:B��ޙ%�[:B:�s�-Qr�M�����ؒ�Y��\ Bƙ��c�l�X˻9�n�cLI��^��Xa)F`m���Tg���yQ�u�����D.(5V�|��.(��=�e��]��|��p�1�ܴyX�
Un3���q�O�.ŗ���H/˒�M~P�)��Tө8B �(w�,V��*+Y�b� ���S��V'�����������9y���ӹ�X��/[�fY�8Կ?��K[h�VP��ֱu��Y3�R�&�3�m�[Fվu�#�r�O�f��?7�X6T�#K<�6�v�^��ښ��y�U�R�z3����%�1T��'�O�)�}�����v>"��#�K�~QU/���8���D�%o�:����O mdXm6o�aV���hbF���A��>�"�dt�Ý�3r|����
~�+��ՈLS��v��u!���.�	��z"y�s�!Ѿ��>,��(�i�O����DXBw�jb<��`%��ɷ2��}a�P
�-�����j>~\���vM���R�^1�k�n��͕�h2oy������t��62O��kܫ�wO�䲪)��.�����^@ʭB�P�=���Wݝ~l�߆�}74��@�o��u�� ޒ>T��b������QJ?���p�B|���UV�>�ϲ�Й����Ǫl���X_�@�N��T��Ul5�`�S���-ˏ�4���&)��fl��q�˹���/�d��k!�i������H��QdN�B"��ԣU�gMx6Ĉ���F�ي�jÍE���X�����A�K��b�I���%>�k��V"y�$�Zb�H�Bk�t�xh���?�V ��ʍ�zr}�������O�=����^S§3ܱ[�ʛ��7,��Z��>n8{SdC��<��G#�����<,A
�7�-���7~�.�o�SE�( <�h���k�������g&�� �G��ү�e���6k�U�h'����&H@4��s�v����XC�74���P���r��\剤u���bu��A����ð�_��/l�����R�ҕM#�Dx;�#\#J!�Y����:�p�1r-EG}��ǂ�%&�������T�r<����� �����s���֛o�Y��{������w1�ۈ.|hc@Nm���"� �C�I�/xX9��6����0���T�6bP@p�c_�꿪s{B�P������x��d��婵��]e�������#�T`�G���w#&V��zHD��\7��Ջ�my z��՜q��o����7�H����LD�MMWڕ�Ln�6��n"�D�?��.7~6v[�s�1�u]��9k:DհJT]�v��̷�ǫ�V�J��$�k���Vx���7� b�o-��Ƴ=�b�j���!�HvH������=�����9m����ST����&�t.Z�G�W �k�����T��8hj�uk��R_H��sH�b�-c���&m���Ǧ�.HK�iE�����'�M������?G��~pZPv��z"��V����ra9O�I$�)쥽+����?y9�a	�5���+�Kq��;Up���C[Z�`+\g@{@�>y�6��L���̗:�WyѪ>�%X��/�g{��8{�v�L�9�@[V��I���*/���<�R�d��TU�@�%�H�$�I��C�'�F[̸@���E��R*XßEۤ�X�G��Oh���>�|��D�'�=��	�y��_�����T��o B~�N���Ӕ�$JѢ�cUg�9 0:�:�|G�it MHۏ�-Y���"�Rq��NK��a3o.�ʬZ��Ly���5 ��RPΉ��w�ʥ]��ֳ�6�Z���H�n!L�#ur�dӚ�&MX؇i�bt�M�΄�Z�/��#nV���p_�2�-MSv6
',��4Ӥ,0Ե�F�� ��FttD�Mt��ӿ�F��/-��a�0���)·E��l3$Bou� 2�!�ʻ�9������(�I_�ަ.����n4�DY�[Pu0t���>��S��d���@�֜�Ef���)�3o;-���@�1���!�Â��5k��K�f<�����1�@�<����LP����ڕ�+����/6L�y �(� D�J��Hl�����3��g�.�o6�5ɯy�5��c�IS��9�
�ō���%��J��[�1�M<�Xf��O��l�[g�߬�<B1�b��6�?���]a����`t��קh�?�r�L�FA�:^�?l�N�\�fT�=��C��L�b���%S�&�����ئ�ϱ�{P��:ph���8+���)���(j|)��hg-��xVG�_}��@�J���l�6�
v���,��p�0.'���c�9�Ggʎ ��n�i��Bf�����D���0�]��d��1�ʴ{��
��A����	�#� �`���>A��H�~�a���%���h~}���/�(���X�/0���9}➷zHj�r�Z߰#B�6)�s��s��w���}-N�$e)��^�u���B��U�|���TK�s�e£3Ǹ�q����YrТ]Z�ے[T>_Rbr��0݅p�H��9���W6����A`� a��D�;����F�7yA-'��!�D����Z�;�������P��I�Vl���J/s��<�S�m�6vk]>z��S�J��T%&�u�0�����o(g� ���(�����n[����7�^N��s�4�00���ȴ��\�3�*2��[󋂛�Kk�ت�m&v�,�,����|`Ǘ��-2} Q����$��e��]�i�PCة�̉k�N��zm;���{1TVd��Ҳ��@{��h���vq��*��*��AX(]K-�+K�=�7�Z���s[HݳN��͒Z��O��~oV��wKT�n�0&]�aA*�;YB5b�F�L��#OPm+�N�+Sn�~96�Z��
�m]��L�j�I�(�;����i��~!WiqN��i�j��w�ohe0�v��Z^�b��GguoCb׽��	q��pȹ��Aڗ,�j$8��z�(��,�:o��Y?����jVڟ:\�>S*cElߣ��͔�ask����x���W5��u7��7r�)21�����h�΄۠G�N�ɗo���Z��l���n��_������)F.懄=�d&�/���e�"w��y�:��^+DA�-	��"o�&�K9_J����9ha��?��e"\����)�ɡ�,���ykn{����jr(��F���c��\�h��E@)��T�T�R� 
B0p�#��#] �=+��v��jZ}��:X�`0�_%8��s��
=#3sUgdG����l������oM��z�h�q0�b�����X�!܌;�M���d �O���4��s���tf�z1�/+��M��%���-�!?�4��*��_3aa���ӿ���8��,��R7����k(c�ӷDX�鄞נyG��(*��@�^)#	����7����ڳ�p�fa՜i�#ꂊ*4�εo�i4� �҇	�W�4&��a4���'��|ٞ�YM�\,p�u�i�a2��K��9�� ��IP����xa���}X�r^Ţ��l�d�w���f�:~"VT:�=�ސ���)m:/
��d��m�n��p����[�::aep�a`|��Z�}���ʒ1���N=Q��S6���ģ�PF�g��2�-���h�C�sXI%P�}G�5A�rCv~�����5��B���Ѱ��e\̰�p�Lˤ�pj�P��?SH�GZD����c'.���h�D����>WK�;�0E��K���h��J�=VQ£b����l���0gg<m����)�G��@���M����;�����?l+}'?8��� J�`#�ԡ�*��C����NbV��ҎU`�&M����"��W0d���Vџr6����`�I�X�}�58�P]�A��"�T�_�T�i���.���m����%�W�ڀ5��Y´A�e7�L~y@,j�-��NX�Gh�!f���g�O}#�O9�!�R)��3�����EY�� b�}�R�T�3&0�A����*���PiH�K��t�
�-�Q��JT����=M� e�J�<�r{F%������,�o2
����Ŧ���B��� v�w5��.u`��b�0�7KZ��{6�$HG���W�j�>��m�.���a����+!լ�����=��	����>W�L+*�]`��I<P���xfRo��H$���Ӝ� ����������&O܌��Ƿ܌�D��S�5{��2,ꃩ+���=^=" �b���F�"���؂V7=����{�����Q7S��
��,��6��.n� �(�ƽT�
U2E$�ٵb��9�U	�]���K����a)�g��S����;�L;�|�c�+��)��3~�؋��>�u�	RPѢ����&����;���|�s�%jX�8�:v1䰭�co�B��H����#S	nܶu9.��ҧ���XYw��D�ixM0�Pٜ�"Ý0�O�gU�o��������Zs�X��T>�f�l��Z��A��-�w!�����c����'�A��+�|�꾂��M��v<ܾ�L���A��u7��w�)<���1����+�q}�G� ؏�>m�5����._�sL����N�;.p�O��h�-x����ځ�E���6g���>�Q�^?;�L�G$ʆ~�i�Z��8`F#x�tM���̂yg�t|~��m�b����k��~u��*����G9����܇M(Y�=p�8�O�Ou��I�B7�D>�z�L�~XI��	��;��S|)����ʷQS/J0Ҝ]�C	2p�>_3�J�:0���~�<t�=���=��O�[%���rq>�v�ڡ"�{�z%�@c��I����]�aWaL��Yte^Hgu�ZͲ0��$ʶ�Ȉ��u���掘�.e�L�c�'�]�I;�)ai�[��ͣŤ�K�v��d�)**�jU��ڔK<��ṣ/��(����Grb��������OL��BOU�B�/�[�H�����{+e�m���u�[Iby���K7��.�Ʋ5F����{��y@&�؉�k$̤3K����gmcgH0T5�8LB��G�179���Ay���)����|�,O6�ŭ!�m9��A��	S���YD��u��fZI2q�� -�z�ƁL�1�r��r�Wc
х���I��f3J�*�%�a�GUG��| q���E7f��Z�M�:2���������G�KH�~+$ˇ���BȮ|�]��B�G�&d*�O\_\8w�Q��I�<:? �R6�V���*�xaQ����/e�C�)\D��3�� �k�ƠtAu��� �G~��;�>τ��v d�����
xY)nN�KEZ��^���]�^�`?�n�s/�P?ݠE)yІ��};T��~���N���� y2}=�}��ӣ��kI1�����uP��ETp��f,xh��g��R��u��ܼѡj��C�p��(��L��&��-#3�#y�ۤ��+s�"�f��s�(r��O_2���jo��]|��2�r�^�[^={���I9��LD�"2o��E�퍪:�Ъ�oFc%�j]��Y��@�P���[iG��s
NREBǾx��ABɞ'����m���^2��m�>o�t�#K�,x	eO��X
��Z�J�Ŏu:m]�% �����0i�T��������Hƫ].JZ)�B>�&m�dۃ�[E��_��.9I����:�(״��|�~��ץ�^;���P,�IИ��u��Y}�;���9�����[�b~��^�o�w�G"x2�rjnd����c5.{#��K|�O8�U�A�&����C7{�]i�����[���d�\�?z4q������>��H����}�li�I���dSw���Q��G2���	����E=eH!�a��
i��e]���R�ċT��M�d|G�� ��#0�NX ���~	D�̓�H� z��T;!���(���� *rs���Hյ׏ru<O`�lM�JB70,~���+�x�Z��2&���(�$lP="�6*;��1i׹U%�ߔo�e��d��o���T��GEN ���ܵ]b"J�I~���dq��/�����ot���E��4�6��je�l�`� �M��c����iD��is��/�o�u���Np₎��:�VMc�V��U���b9-��mMn�9����m{�� "+�Xu����2�\s��F��aRm���xY��bN
K�!(���xL�E�� -K��Y����3�wO���a���eiā�)�%�}��-߿]ؠ��a[͇B�z/j�Lؖ��2K>dN��̃��z����Ҷ;c��d;�w6/{��47}�0,�Y�X(� 
�pq,��3"�)�Up�HH��� A�G������ؾn���Z�	�������]e�V>svB���!�5�K|^�B0�S&@�)ba�U��M��^���<�����N\�A?�c�0�1˚�Q?��슿7�q5MeF���GI�͎�w�>��6�j�*X����� ��1��Jq1Z�ꄁ+��>e�ޅ�n"T�k;mYjP����U'7A�c_eq�"u�c�!	��v��枝Ŗك_(�N�ߎ�ѧ�bi�.˘�����\uȝ����Db���Oj�S�����!,O�v_W�r3;�gcS`�}#�������3,:�s���smϕwb�9$.�`j*��z���y�L��g5_>�����5!��Ƅ���`��R�E�g-�zb�e�[]�=5�0�R�M����~�����q��/|�h��e���Xoc���Gю�c���Y����W���{w�0K3��QW�!��?1�xF�x���1E�]�ؿ4�6K��ydjLO�U�����I:d]w
Bfy���X7��;����]�&#�mV:�?�uFG<43ʞ*��!���}�4��5��E�(!�6��)�(��H$��\�U,�SND #�+mʂ*%^�Za��0�]��]��^�G�}k'+�v��8S�P�-�J��a��Ys7��Ѵ��:>�2��.��3
�ر�f���_������d���4�Xu�~������66�O��O���4��+��8���C�Ik��BO����z����x�0���Ƶ$�+08�o0nGZԃ�j�OF�N�|4Y��#�&��������M��?R|Q����d�)��Zea�;�w�>m坸�'���<O&B��7M�	��ۭ�°=�Ϥ`�`�u��m�>Zu�dc��£dQ��>�����0�Y1�����_-N�}uC�-����TQf1�Hl����u>��W�Ӷ�&G�8pv࿞�<I������7��8��
u7$�d����=ڣ�k?�R�-���+���CF~o�}Z�����-V���=��p^x
!��Y|� \����'F�u#g�ff�/�v�^6N��	r��I7���Nk ����qP��w��͉<g�<=�ŝN�X��n�����e��_���&���Am�. �qBfH5<k���O��}*�mu�Fǰ}M���m_��Pcփ�}��W@c�|�W��Ǿ����]�|��i������y,��q��F��r�s���ч	��:
�^���LBsث�_S�=��4h�&C8���Z`@ GG���Z7r��\�k�.P����Iݕ��.:@���������.�{����㲰�U_����~^�o��eܝ�� ��
z�/.���^��r���F�	P��.B�9Tv�}�ͥ~w%Rɣg�U[kxE��lM<�����[i)]��.�D]��Qih@��ܼ����*Sj��e|��M�����;�Y�W�=��_��k
ä���(�j`�����1(6u�<8ۋ۸Gͣ�.!Y���=����S��!�?��ѧ�-��l?�w�Ї��3�C��J�� 4�i�~z9g��+��R�p���x�i�Қ\� ��q�Xd��p8y�<Q���g��@hT�P�}y��䌱����k��H1���@~�´e�漮��%��3,0&�;k��WKN�Em��:���o�x-��4��?��=�_�m\�k2v���9��Y�o$�(����v�-9�sf/����e���4b�,"r<�N�A�䘹��nW\�g�,����]ӔU�υLr�Ie2�V6�xa���F���Ŀ�Q�UH�ELgLU��n�%�.��f��q>%젭�is)S��k�����!sli���~.&���j�L�� h�MOT�@h{���g���iF������`��śր>����D�*|	�%a"޿��RUC�͚A��9k����d�zc��G�`�0GȒ�w���~���I�]3R�ۓ[�FD�T�c�t��枸���߿��֍D��6�oZ��7T�G-9���fa�d�O(�k�_d�.����k��R0A��a�!�6����Փu����gЙ$�9p��8��q�h1�������9��x��w��Z�YaG/#��|����
�#w L�̻#�yл5n��!~��,�O~��kc�aϟ�p)��F�<��a;;e2s�q��3��W����X��a {��� 11l �E�� ��l�]��"\	�
�*3M�'"-�CPy+;_D&<�D;#�BYH�r:<K����#2 ��;������L�2��'T>>6����VKA�_2C��>�"�/�E�����p���DY�7�>3�t�S��~�i����c&�Ta~��?�ܯh��\� �1�:����2l4�fݖ��U��L�W⁄��RD�R(����s�93��|.2X�!cn�ݠ��l��fE�-yk?�y��$�'��8%k��l��p�Ӌ��9>� �)2�`��^�w�eB��6��Ʉ`S#uk����f��H��q=3I�����ډg :y�AƧ�<"���x&�� Ts�7z�dS��j2P�@�|H����_��˔��� �3 OL���R�n߃D���Z���b�3T�N�9R|�0�ːg�ջ�YTD���>�^�ÁՇ�e�g��K#^g�N���^�z�R�%��ə�h�r����qT�#BMqLl���� �ٷ����s�g>QpjOU�g_������S&>�$]�����D�\a�=����RhBx��m$�ZP�(vȏW�I2���kG��J���=�p������r@9���М-H�#{z`	�.�,�b�~T���\�,?��VjI��e��
6�.��a"�wN�L�s�I�����	�F!Rzˊ�,�P�/�e�
��~��@8�~G�f�淠�V��Җ������)?=���䉾�.�]�����+�X㝌���
���Ą�DU�u�6xO�k��T�Ò�
��c��N)@�戒���!Cm��ej&�Rs�;�6*���k�"5��_o��3W��/l�@e	��hP<��DK�AL hNu{Ϋ�^��@a�fV��kĢ?2G\ܨV;�>^��ypȲ}Wđ`���I��z��o�>q<&�m����8@�N�lq܌��L���r�5�S#��