	component cpu is
		port (
			buttons_export                             : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			clk_clk                                    : in    std_logic                     := 'X';             -- clk
			hexes_export                               : out   std_logic_vector(27 downto 0);                    -- export
			hps_io_hps_io_emac1_inst_TX_CLK            : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_hps_io_emac1_inst_TXD0              : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_hps_io_emac1_inst_TXD1              : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_hps_io_emac1_inst_TXD2              : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_hps_io_emac1_inst_TXD3              : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_hps_io_emac1_inst_RXD0              : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_hps_io_emac1_inst_MDIO              : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_hps_io_emac1_inst_MDC               : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_hps_io_emac1_inst_RX_CTL            : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_hps_io_emac1_inst_TX_CTL            : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_hps_io_emac1_inst_RX_CLK            : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_hps_io_emac1_inst_RXD1              : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_hps_io_emac1_inst_RXD2              : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_hps_io_emac1_inst_RXD3              : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_hps_io_qspi_inst_IO0                : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO0
			hps_io_hps_io_qspi_inst_IO1                : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO1
			hps_io_hps_io_qspi_inst_IO2                : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO2
			hps_io_hps_io_qspi_inst_IO3                : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO3
			hps_io_hps_io_qspi_inst_SS0                : out   std_logic;                                        -- hps_io_qspi_inst_SS0
			hps_io_hps_io_qspi_inst_CLK                : out   std_logic;                                        -- hps_io_qspi_inst_CLK
			hps_io_hps_io_sdio_inst_CMD                : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_hps_io_sdio_inst_D0                 : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_hps_io_sdio_inst_D1                 : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_hps_io_sdio_inst_CLK                : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_hps_io_sdio_inst_D2                 : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_hps_io_sdio_inst_D3                 : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_hps_io_usb1_inst_D0                 : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_hps_io_usb1_inst_D1                 : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_hps_io_usb1_inst_D2                 : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_hps_io_usb1_inst_D3                 : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_hps_io_usb1_inst_D4                 : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_hps_io_usb1_inst_D5                 : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_hps_io_usb1_inst_D6                 : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_hps_io_usb1_inst_D7                 : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_hps_io_usb1_inst_CLK                : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_hps_io_usb1_inst_STP                : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_hps_io_usb1_inst_DIR                : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_hps_io_usb1_inst_NXT                : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_hps_io_spim1_inst_CLK               : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_hps_io_spim1_inst_MOSI              : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_hps_io_spim1_inst_MISO              : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_hps_io_spim1_inst_SS0               : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_hps_io_uart0_inst_RX                : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_hps_io_uart0_inst_TX                : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_hps_io_i2c0_inst_SDA                : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_hps_io_i2c0_inst_SCL                : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_hps_io_i2c1_inst_SDA                : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_hps_io_i2c1_inst_SCL                : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_hps_io_gpio_inst_GPIO09             : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_hps_io_gpio_inst_GPIO35             : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_hps_io_gpio_inst_GPIO40             : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_hps_io_gpio_inst_GPIO41             : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO41
			hps_io_hps_io_gpio_inst_GPIO48             : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_hps_io_gpio_inst_GPIO53             : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_hps_io_gpio_inst_GPIO54             : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_hps_io_gpio_inst_GPIO61             : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			img_cpu_reader_0_cpu_rdy_cpu_rdy           : out   std_logic;                                        -- cpu_rdy
			img_cpu_reader_0_get_next_pix_get_next_pix : out   std_logic;                                        -- get_next_pix
			img_cpu_reader_0_img_done_img_done         : in    std_logic                     := 'X';             -- img_done
			img_cpu_reader_0_out_state_out_state       : out   std_logic_vector(3 downto 0);                     -- out_state
			img_cpu_reader_0_pix_rdy_pix_rdy           : in    std_logic                     := 'X';             -- pix_rdy
			img_cpu_reader_0_pix_rdy_out_pix_rdy_out   : out   std_logic_vector(31 downto 0);                    -- pix_rdy_out
			img_cpu_reader_0_pix_rgb_out_pix_rgb_out   : out   std_logic_vector(23 downto 0);                    -- pix_rgb_out
			img_cpu_reader_0_pixel_data_pixel_data     : in    std_logic_vector(23 downto 0) := (others => 'X'); -- pixel_data
			memory_mem_a                               : out   std_logic_vector(14 downto 0);                    -- mem_a
			memory_mem_ba                              : out   std_logic_vector(2 downto 0);                     -- mem_ba
			memory_mem_ck                              : out   std_logic;                                        -- mem_ck
			memory_mem_ck_n                            : out   std_logic;                                        -- mem_ck_n
			memory_mem_cke                             : out   std_logic;                                        -- mem_cke
			memory_mem_cs_n                            : out   std_logic;                                        -- mem_cs_n
			memory_mem_ras_n                           : out   std_logic;                                        -- mem_ras_n
			memory_mem_cas_n                           : out   std_logic;                                        -- mem_cas_n
			memory_mem_we_n                            : out   std_logic;                                        -- mem_we_n
			memory_mem_reset_n                         : out   std_logic;                                        -- mem_reset_n
			memory_mem_dq                              : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			memory_mem_dqs                             : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			memory_mem_dqs_n                           : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			memory_mem_odt                             : out   std_logic;                                        -- mem_odt
			memory_mem_dm                              : out   std_logic_vector(3 downto 0);                     -- mem_dm
			memory_oct_rzqin                           : in    std_logic                     := 'X';             -- oct_rzqin
			reset_reset                                : in    std_logic                     := 'X';             -- reset
			sdram_addr                                 : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_ba                                   : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_cas_n                                : out   std_logic;                                        -- cas_n
			sdram_cke                                  : out   std_logic;                                        -- cke
			sdram_cs_n                                 : out   std_logic;                                        -- cs_n
			sdram_dq                                   : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_dqm                                  : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_ras_n                                : out   std_logic;                                        -- ras_n
			sdram_we_n                                 : out   std_logic;                                        -- we_n
			sdram_clk_clk                              : out   std_logic;                                        -- clk
			switches_export                            : in    std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			touch_uart_RXD                             : in    std_logic                     := 'X';             -- RXD
			touch_uart_TXD                             : out   std_logic;                                        -- TXD
			vga_CLK                                    : out   std_logic;                                        -- CLK
			vga_HS                                     : out   std_logic;                                        -- HS
			vga_VS                                     : out   std_logic;                                        -- VS
			vga_BLANK                                  : out   std_logic;                                        -- BLANK
			vga_SYNC                                   : out   std_logic;                                        -- SYNC
			vga_R                                      : out   std_logic_vector(7 downto 0);                     -- R
			vga_G                                      : out   std_logic_vector(7 downto 0);                     -- G
			vga_B                                      : out   std_logic_vector(7 downto 0)                      -- B
		);
	end component cpu;

	u0 : component cpu
		port map (
			buttons_export                             => CONNECTED_TO_buttons_export,                             --                       buttons.export
			clk_clk                                    => CONNECTED_TO_clk_clk,                                    --                           clk.clk
			hexes_export                               => CONNECTED_TO_hexes_export,                               --                         hexes.export
			hps_io_hps_io_emac1_inst_TX_CLK            => CONNECTED_TO_hps_io_hps_io_emac1_inst_TX_CLK,            --                        hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_hps_io_emac1_inst_TXD0              => CONNECTED_TO_hps_io_hps_io_emac1_inst_TXD0,              --                              .hps_io_emac1_inst_TXD0
			hps_io_hps_io_emac1_inst_TXD1              => CONNECTED_TO_hps_io_hps_io_emac1_inst_TXD1,              --                              .hps_io_emac1_inst_TXD1
			hps_io_hps_io_emac1_inst_TXD2              => CONNECTED_TO_hps_io_hps_io_emac1_inst_TXD2,              --                              .hps_io_emac1_inst_TXD2
			hps_io_hps_io_emac1_inst_TXD3              => CONNECTED_TO_hps_io_hps_io_emac1_inst_TXD3,              --                              .hps_io_emac1_inst_TXD3
			hps_io_hps_io_emac1_inst_RXD0              => CONNECTED_TO_hps_io_hps_io_emac1_inst_RXD0,              --                              .hps_io_emac1_inst_RXD0
			hps_io_hps_io_emac1_inst_MDIO              => CONNECTED_TO_hps_io_hps_io_emac1_inst_MDIO,              --                              .hps_io_emac1_inst_MDIO
			hps_io_hps_io_emac1_inst_MDC               => CONNECTED_TO_hps_io_hps_io_emac1_inst_MDC,               --                              .hps_io_emac1_inst_MDC
			hps_io_hps_io_emac1_inst_RX_CTL            => CONNECTED_TO_hps_io_hps_io_emac1_inst_RX_CTL,            --                              .hps_io_emac1_inst_RX_CTL
			hps_io_hps_io_emac1_inst_TX_CTL            => CONNECTED_TO_hps_io_hps_io_emac1_inst_TX_CTL,            --                              .hps_io_emac1_inst_TX_CTL
			hps_io_hps_io_emac1_inst_RX_CLK            => CONNECTED_TO_hps_io_hps_io_emac1_inst_RX_CLK,            --                              .hps_io_emac1_inst_RX_CLK
			hps_io_hps_io_emac1_inst_RXD1              => CONNECTED_TO_hps_io_hps_io_emac1_inst_RXD1,              --                              .hps_io_emac1_inst_RXD1
			hps_io_hps_io_emac1_inst_RXD2              => CONNECTED_TO_hps_io_hps_io_emac1_inst_RXD2,              --                              .hps_io_emac1_inst_RXD2
			hps_io_hps_io_emac1_inst_RXD3              => CONNECTED_TO_hps_io_hps_io_emac1_inst_RXD3,              --                              .hps_io_emac1_inst_RXD3
			hps_io_hps_io_qspi_inst_IO0                => CONNECTED_TO_hps_io_hps_io_qspi_inst_IO0,                --                              .hps_io_qspi_inst_IO0
			hps_io_hps_io_qspi_inst_IO1                => CONNECTED_TO_hps_io_hps_io_qspi_inst_IO1,                --                              .hps_io_qspi_inst_IO1
			hps_io_hps_io_qspi_inst_IO2                => CONNECTED_TO_hps_io_hps_io_qspi_inst_IO2,                --                              .hps_io_qspi_inst_IO2
			hps_io_hps_io_qspi_inst_IO3                => CONNECTED_TO_hps_io_hps_io_qspi_inst_IO3,                --                              .hps_io_qspi_inst_IO3
			hps_io_hps_io_qspi_inst_SS0                => CONNECTED_TO_hps_io_hps_io_qspi_inst_SS0,                --                              .hps_io_qspi_inst_SS0
			hps_io_hps_io_qspi_inst_CLK                => CONNECTED_TO_hps_io_hps_io_qspi_inst_CLK,                --                              .hps_io_qspi_inst_CLK
			hps_io_hps_io_sdio_inst_CMD                => CONNECTED_TO_hps_io_hps_io_sdio_inst_CMD,                --                              .hps_io_sdio_inst_CMD
			hps_io_hps_io_sdio_inst_D0                 => CONNECTED_TO_hps_io_hps_io_sdio_inst_D0,                 --                              .hps_io_sdio_inst_D0
			hps_io_hps_io_sdio_inst_D1                 => CONNECTED_TO_hps_io_hps_io_sdio_inst_D1,                 --                              .hps_io_sdio_inst_D1
			hps_io_hps_io_sdio_inst_CLK                => CONNECTED_TO_hps_io_hps_io_sdio_inst_CLK,                --                              .hps_io_sdio_inst_CLK
			hps_io_hps_io_sdio_inst_D2                 => CONNECTED_TO_hps_io_hps_io_sdio_inst_D2,                 --                              .hps_io_sdio_inst_D2
			hps_io_hps_io_sdio_inst_D3                 => CONNECTED_TO_hps_io_hps_io_sdio_inst_D3,                 --                              .hps_io_sdio_inst_D3
			hps_io_hps_io_usb1_inst_D0                 => CONNECTED_TO_hps_io_hps_io_usb1_inst_D0,                 --                              .hps_io_usb1_inst_D0
			hps_io_hps_io_usb1_inst_D1                 => CONNECTED_TO_hps_io_hps_io_usb1_inst_D1,                 --                              .hps_io_usb1_inst_D1
			hps_io_hps_io_usb1_inst_D2                 => CONNECTED_TO_hps_io_hps_io_usb1_inst_D2,                 --                              .hps_io_usb1_inst_D2
			hps_io_hps_io_usb1_inst_D3                 => CONNECTED_TO_hps_io_hps_io_usb1_inst_D3,                 --                              .hps_io_usb1_inst_D3
			hps_io_hps_io_usb1_inst_D4                 => CONNECTED_TO_hps_io_hps_io_usb1_inst_D4,                 --                              .hps_io_usb1_inst_D4
			hps_io_hps_io_usb1_inst_D5                 => CONNECTED_TO_hps_io_hps_io_usb1_inst_D5,                 --                              .hps_io_usb1_inst_D5
			hps_io_hps_io_usb1_inst_D6                 => CONNECTED_TO_hps_io_hps_io_usb1_inst_D6,                 --                              .hps_io_usb1_inst_D6
			hps_io_hps_io_usb1_inst_D7                 => CONNECTED_TO_hps_io_hps_io_usb1_inst_D7,                 --                              .hps_io_usb1_inst_D7
			hps_io_hps_io_usb1_inst_CLK                => CONNECTED_TO_hps_io_hps_io_usb1_inst_CLK,                --                              .hps_io_usb1_inst_CLK
			hps_io_hps_io_usb1_inst_STP                => CONNECTED_TO_hps_io_hps_io_usb1_inst_STP,                --                              .hps_io_usb1_inst_STP
			hps_io_hps_io_usb1_inst_DIR                => CONNECTED_TO_hps_io_hps_io_usb1_inst_DIR,                --                              .hps_io_usb1_inst_DIR
			hps_io_hps_io_usb1_inst_NXT                => CONNECTED_TO_hps_io_hps_io_usb1_inst_NXT,                --                              .hps_io_usb1_inst_NXT
			hps_io_hps_io_spim1_inst_CLK               => CONNECTED_TO_hps_io_hps_io_spim1_inst_CLK,               --                              .hps_io_spim1_inst_CLK
			hps_io_hps_io_spim1_inst_MOSI              => CONNECTED_TO_hps_io_hps_io_spim1_inst_MOSI,              --                              .hps_io_spim1_inst_MOSI
			hps_io_hps_io_spim1_inst_MISO              => CONNECTED_TO_hps_io_hps_io_spim1_inst_MISO,              --                              .hps_io_spim1_inst_MISO
			hps_io_hps_io_spim1_inst_SS0               => CONNECTED_TO_hps_io_hps_io_spim1_inst_SS0,               --                              .hps_io_spim1_inst_SS0
			hps_io_hps_io_uart0_inst_RX                => CONNECTED_TO_hps_io_hps_io_uart0_inst_RX,                --                              .hps_io_uart0_inst_RX
			hps_io_hps_io_uart0_inst_TX                => CONNECTED_TO_hps_io_hps_io_uart0_inst_TX,                --                              .hps_io_uart0_inst_TX
			hps_io_hps_io_i2c0_inst_SDA                => CONNECTED_TO_hps_io_hps_io_i2c0_inst_SDA,                --                              .hps_io_i2c0_inst_SDA
			hps_io_hps_io_i2c0_inst_SCL                => CONNECTED_TO_hps_io_hps_io_i2c0_inst_SCL,                --                              .hps_io_i2c0_inst_SCL
			hps_io_hps_io_i2c1_inst_SDA                => CONNECTED_TO_hps_io_hps_io_i2c1_inst_SDA,                --                              .hps_io_i2c1_inst_SDA
			hps_io_hps_io_i2c1_inst_SCL                => CONNECTED_TO_hps_io_hps_io_i2c1_inst_SCL,                --                              .hps_io_i2c1_inst_SCL
			hps_io_hps_io_gpio_inst_GPIO09             => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO09,             --                              .hps_io_gpio_inst_GPIO09
			hps_io_hps_io_gpio_inst_GPIO35             => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO35,             --                              .hps_io_gpio_inst_GPIO35
			hps_io_hps_io_gpio_inst_GPIO40             => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO40,             --                              .hps_io_gpio_inst_GPIO40
			hps_io_hps_io_gpio_inst_GPIO41             => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO41,             --                              .hps_io_gpio_inst_GPIO41
			hps_io_hps_io_gpio_inst_GPIO48             => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO48,             --                              .hps_io_gpio_inst_GPIO48
			hps_io_hps_io_gpio_inst_GPIO53             => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO53,             --                              .hps_io_gpio_inst_GPIO53
			hps_io_hps_io_gpio_inst_GPIO54             => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO54,             --                              .hps_io_gpio_inst_GPIO54
			hps_io_hps_io_gpio_inst_GPIO61             => CONNECTED_TO_hps_io_hps_io_gpio_inst_GPIO61,             --                              .hps_io_gpio_inst_GPIO61
			img_cpu_reader_0_cpu_rdy_cpu_rdy           => CONNECTED_TO_img_cpu_reader_0_cpu_rdy_cpu_rdy,           --      img_cpu_reader_0_cpu_rdy.cpu_rdy
			img_cpu_reader_0_get_next_pix_get_next_pix => CONNECTED_TO_img_cpu_reader_0_get_next_pix_get_next_pix, -- img_cpu_reader_0_get_next_pix.get_next_pix
			img_cpu_reader_0_img_done_img_done         => CONNECTED_TO_img_cpu_reader_0_img_done_img_done,         --     img_cpu_reader_0_img_done.img_done
			img_cpu_reader_0_out_state_out_state       => CONNECTED_TO_img_cpu_reader_0_out_state_out_state,       --    img_cpu_reader_0_out_state.out_state
			img_cpu_reader_0_pix_rdy_pix_rdy           => CONNECTED_TO_img_cpu_reader_0_pix_rdy_pix_rdy,           --      img_cpu_reader_0_pix_rdy.pix_rdy
			img_cpu_reader_0_pix_rdy_out_pix_rdy_out   => CONNECTED_TO_img_cpu_reader_0_pix_rdy_out_pix_rdy_out,   --  img_cpu_reader_0_pix_rdy_out.pix_rdy_out
			img_cpu_reader_0_pix_rgb_out_pix_rgb_out   => CONNECTED_TO_img_cpu_reader_0_pix_rgb_out_pix_rgb_out,   --  img_cpu_reader_0_pix_rgb_out.pix_rgb_out
			img_cpu_reader_0_pixel_data_pixel_data     => CONNECTED_TO_img_cpu_reader_0_pixel_data_pixel_data,     --   img_cpu_reader_0_pixel_data.pixel_data
			memory_mem_a                               => CONNECTED_TO_memory_mem_a,                               --                        memory.mem_a
			memory_mem_ba                              => CONNECTED_TO_memory_mem_ba,                              --                              .mem_ba
			memory_mem_ck                              => CONNECTED_TO_memory_mem_ck,                              --                              .mem_ck
			memory_mem_ck_n                            => CONNECTED_TO_memory_mem_ck_n,                            --                              .mem_ck_n
			memory_mem_cke                             => CONNECTED_TO_memory_mem_cke,                             --                              .mem_cke
			memory_mem_cs_n                            => CONNECTED_TO_memory_mem_cs_n,                            --                              .mem_cs_n
			memory_mem_ras_n                           => CONNECTED_TO_memory_mem_ras_n,                           --                              .mem_ras_n
			memory_mem_cas_n                           => CONNECTED_TO_memory_mem_cas_n,                           --                              .mem_cas_n
			memory_mem_we_n                            => CONNECTED_TO_memory_mem_we_n,                            --                              .mem_we_n
			memory_mem_reset_n                         => CONNECTED_TO_memory_mem_reset_n,                         --                              .mem_reset_n
			memory_mem_dq                              => CONNECTED_TO_memory_mem_dq,                              --                              .mem_dq
			memory_mem_dqs                             => CONNECTED_TO_memory_mem_dqs,                             --                              .mem_dqs
			memory_mem_dqs_n                           => CONNECTED_TO_memory_mem_dqs_n,                           --                              .mem_dqs_n
			memory_mem_odt                             => CONNECTED_TO_memory_mem_odt,                             --                              .mem_odt
			memory_mem_dm                              => CONNECTED_TO_memory_mem_dm,                              --                              .mem_dm
			memory_oct_rzqin                           => CONNECTED_TO_memory_oct_rzqin,                           --                              .oct_rzqin
			reset_reset                                => CONNECTED_TO_reset_reset,                                --                         reset.reset
			sdram_addr                                 => CONNECTED_TO_sdram_addr,                                 --                         sdram.addr
			sdram_ba                                   => CONNECTED_TO_sdram_ba,                                   --                              .ba
			sdram_cas_n                                => CONNECTED_TO_sdram_cas_n,                                --                              .cas_n
			sdram_cke                                  => CONNECTED_TO_sdram_cke,                                  --                              .cke
			sdram_cs_n                                 => CONNECTED_TO_sdram_cs_n,                                 --                              .cs_n
			sdram_dq                                   => CONNECTED_TO_sdram_dq,                                   --                              .dq
			sdram_dqm                                  => CONNECTED_TO_sdram_dqm,                                  --                              .dqm
			sdram_ras_n                                => CONNECTED_TO_sdram_ras_n,                                --                              .ras_n
			sdram_we_n                                 => CONNECTED_TO_sdram_we_n,                                 --                              .we_n
			sdram_clk_clk                              => CONNECTED_TO_sdram_clk_clk,                              --                     sdram_clk.clk
			switches_export                            => CONNECTED_TO_switches_export,                            --                      switches.export
			touch_uart_RXD                             => CONNECTED_TO_touch_uart_RXD,                             --                    touch_uart.RXD
			touch_uart_TXD                             => CONNECTED_TO_touch_uart_TXD,                             --                              .TXD
			vga_CLK                                    => CONNECTED_TO_vga_CLK,                                    --                           vga.CLK
			vga_HS                                     => CONNECTED_TO_vga_HS,                                     --                              .HS
			vga_VS                                     => CONNECTED_TO_vga_VS,                                     --                              .VS
			vga_BLANK                                  => CONNECTED_TO_vga_BLANK,                                  --                              .BLANK
			vga_SYNC                                   => CONNECTED_TO_vga_SYNC,                                   --                              .SYNC
			vga_R                                      => CONNECTED_TO_vga_R,                                      --                              .R
			vga_G                                      => CONNECTED_TO_vga_G,                                      --                              .G
			vga_B                                      => CONNECTED_TO_vga_B                                       --                              .B
		);

