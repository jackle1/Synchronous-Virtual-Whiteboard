��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3�[�����Pٵ&�����''�qe�-�?
�%w$�W��[��m�w�xH�O�I�	�@����[oVʭM�A��t��B�gx�K���8C��G#h�̾cZ���8���L1�}�L�RZ��L/��W�p���;lB��*�Y��4�%]�Y�:�b�\Yv_f��!P�{
2G�-�Pi���xhB�ё�&���7`��G%����U�^�9���t�M� ���X3���#���u�鉾μr|Wh��h��Kɟ������cG:��9J>:���ϔ"��nE��2�����>pS4s��	�(G4{(S�L�:U�.@�|R0�L8������j��IB�"���N������ys��ė/,ҊN	q�v�Z��\R�w�0xtʎ5x5�������v�7\M�k���%n;c-<�<;�`.���B1�7���[�D�\�A��fIj�)����懋�f�7	�����A�*��k-e%�P��Ҿ��Z�O����K��Qw�K3�\�qRp�2"�Z����&OB�+�s�(�X�q.
��W�W~��'a/Q�k��h�ud����e}j%��tІr�)�j*�(>z�
�+S߶��n���]5��]�����~ L��%���5��V���*Ёg]l�~ˎ[�n�S�S�B����i���Rk�:�QGh"]��UggB�Mc�\��lR]�8����x 7FI5�b���$���㴴Y���CA�SЃz7f�yz�ĺz	Ӡ*���|^y�p��'���!`^��ke%�Q��^��Pٚi6�*�F^9���s���:R8��e�&/�(E���,��Ã�r3KD��>���Q��� ���g�(ǎ��{ibto���b��%H�#h����'�]�*B�_��5������^kX�]~ɣ�A2����FPsm�D�u��-��_��?m�0�;��rN"�D���v�1���\s���y"��ݻ����jk%˺��L�qMۇ�мk�Z�3��o��IE��Z��������)��&�M���3�J�|^��ks��҈�&���gq��'#/�>E�ß3A2�?{�� Z�������K�rHȋ0^�픢�;��C�yH��ű�� X�&ж��A�H���v\ ��G��^p�������"�H0	+D9�}��Q2�4>e_D!T����gE��ؙ�0��Պ�z�<��aF��ܢAF���S�^ĝCw��n���9�>�2��k�0f_ŵ�c�J=�z��Xꭃ�7��i��ϋ�U�Qc��ֹE�%���V۵v�#ޢ�6�� �J'֠"��od<GX�Q�:]*&��+�S���`�?
��o�.x�$Sʽ�#��*��������F�j��~◡�q�?m�I+�Kз��SiDؚ�>�v�C>�%����/,�����3'���������E����`=Q��[���)�F�ìq�4:���1�������6���e�x�RfL���R���p�Y b�x��Չ��4FpS�Y�,a����X�~�cތ��8,�&T࿠�@	3I�pЧ߶���t.�:�xp��3�G��:/��>�T:�A�oLYi���V0�z�5�F,lj���"�c��f1�
l�f)��LSJ}�L��d�XD1Z?�'`�U��֟�2.m���J�Z���y��٫��H�!C�ߘ��w`1i��յf����n��M����d��uɲ���+p��_���ӫ�8pz�b������1�@ǥ�4��՟�R3'#	Y�+�pcU�d�����b��;o���+�Y�D*)�A��~ǌ3��������wV(S�SZ1@
 �w���;w�HT���k� �c��Ǵ�K!O���]�"�m{�R�qϮj�Yg@ �5X�����?�BO�����|Z[d���9�$*(��]�^o�yOgr�%��2�<�ؒ���P���{J^f0���ص�-�a��y_�>��XP��vH�=�N&ä;%�n�q� �qH��$��n�T��YJ�F:H�ʥ�FFU�٣d/-�O]�|�G�P��i��\2,f��ܤH=�m=�0g��}tusy���u7�3r�f��uR쨟���T���V�@!n]� �q�$��ԙ�����}�X���O�41��K6����&:,�P�𔂸CP��U��!���Ʉ�z]{F��釛CG2fH������t?{���3�O��8�Q�r��$[�	c��]Gټ2�m��ty����㢦�P�B���._�G�u�Y	���Ǩ]��E�j��:�(��|���t�8fiv�q����dc�N��y�d�o��������oK�.L-=f=����4\���D����| w�%�p�9G��s��.�}�Cm����ndv8��9&������Gl�[����	�/���=	��~���*���R1�F6HI�v�mo��&��P��u�IF�-�ȶԘ��)ɷ�1W��F=?�r�pD�^2fS�J$��1�Q0��x�#M�W������6o���t,�g\� ?+8�YJ������W
�&r���]��S���b>a_.�p>���c����	��_�v>�`Z����y��"Y�hx��v��XBH|���nl���Z�J`u�頂6s�cy�	d�'�x�,K��-g-���[(_o<K�+�t��.�"ě�Ѹ���z^;���*�4R��馜G���U#.��g���+L�|z>��α8�<;±���L�����D�1ˢ33��w��X�r��.pŪ���ܜ@��!�{G�M� �8�t�]g�x��z��r�JʜQͷ=kJ�tc��o�8�v��W�%jN貍c���q.1x"���Ȁ�ND��rq�(�j�Y�MF��7ϩ؄�ëF[�����{O��7FA(/�#:�ާ��<�dVg�,-|& �}a��1D!��tlX��ѢP#�s�<�b����p�T��܉׷w6�>��ͪ���䴗5m���:Q�_��Vv��O�s�@�Ċ�:�u��"��Ͼ�x�Ģ�R����� �M1��`�Ŀl{�H�G�3e��R�5y\��{7�Hg�o�L�Q��_M#�Gwy� 厮�����d���0s�\�	ά��ޤ_�����7*`o@r�4�_��O�m�ۄ<�&��N��Yjc����=mHA�E/���6��[��p�Ǻ�6�Жr�d�՚2�i���\I̒r��̾��y��K�7�Bi5��Q�
,�7�#��pu^��BU��:{���0>����y��W������3O�Ǜ����(_"����ɝ�B,_(?��������2`��u�3�}l�X��b!3�n�����]d�)�n+�|Շ@ۨm V�j?�a�Nb�	㰹}�C4��Gw˛$�Z5bE��R�����+6���%:8\C��m'#T�rZo�e��p�ݕ��mJ<�HP��M�\���5Q+�{e�n�<Y��$�M�bG�D�f�������H��T��J��o0?��_�E0��?Pvq��+� ��j�22fPL�*%>n��VQT� ew�4����贇�\ES��ݽ,�@5�i��%u
e����4gg���)�\ ���C��4'ÁZ����C
L9n|,{��,��%������/-� LȶڗUm�yT��ʹ]�Aup��i�uzeW=��;{�w��%T�
\bk}����~&��<�~��yiZ��U�0Ӕ�	�bַ��`F�8���x�n�!��k[kn[�����SP��:���edH�V�R�|��(������c�$U���|J�����1����b�8�8��Ow&���S%���d>�9�|�-����~(ӈ��k�e�}~2�4�` �I���g�����+�|I�LuFgb��\X��W仠�G����B��@�,�}Py�u��VT��܅7�|�XKa]L�3����L�V�@F�p� c���*u v��O�
�Rn��=^#jh��t���\v��z[(��I�Y�z�z9<ύ���q>,^�jeU{�gf�_��$��e�>'{O�bM
���1�����9/	����b��̳S��8�J����U��j��z���Pp<#�-��Ǵus��v:y �9c�O�_���G�����qߋM��&N]�>��Dq�ݑ����|Bj�	�J&�֞	� W��{X�ͼW���s�\�a���*�v,�1-��ʉT<�*K��!ϊѴ�9�d�� ����*�q.�*ei7�w��U�dh"T��P�KP�� ��i ���=���49�H��O�%�����L�-�c�4��"O=X�����G�"�����Kk�#X��bF�1	��16E�A�9��n���D�P�_�����0���VO���~ې����,����ĉ�#��w�9[�!Ʉ8�k���q���؁|S�t��by�"ϰ8��گG�i�ŷ���w�ޚ > �f��m�d�S�ʜ�՘���Ro��./�׬ŷ�c}>%h�z�I����'�ᇑ�'�`���{ٜ�S&vT������]�{+�a9fwz�M��V*X�Hw`.���K��?�a�(�zirJ(�1��O\X�;�w�a���1t�+���N2�>���MXH��k�\?�%���y����͞P/�npyN�8���Lw]�����/4�v �����Zc�F=I����F�0���d?�tMz�ܡ�m!�����8�}�IĿ���(�������{h���{��s9$H�n5sR���GA��CPy�����c��A���D7�1c^@n+�߉>����5�D��r�'lO6��Gt�u���[ �4�U�9`�o{�O�p����C?��L��H�p]V*�8d\�<��t���ލ�`�ώ�����~0,�Ξ�͏W��8O\鵦�t�-nmU�m�D��k)�Z�t|��k4��GLb9SZ?���%)tg�$�X������p̟�G}B_lk+�(�9>7��	������:���������%h�#��^ �A�e�̟���+����@���}�]k+���=�O� A�iG��־!�ȋ^(r�@骸��������������}�@�`1:s��g�>�U�d-���ؚt(ɒ��p�� +D3@j����� �ʖ��d1����'C6]*�����[Ne5D���[
��	hy��v����Q��+���\�W�+�	1����!��(�I�w&m�p#����!ięcB��f0�_	�be˷?�Ƴe�q1�4�	WT���s�YS<D�ɴ�������x8JT.��h�A ��!�s�	4t#��:��S�һ�N�tM�.�u�(����+fֶ���|�+J��ϧ�q�&PtW�����O�W�H7�������&����Py�����y�#�f?8����? ���eh�,,�
�$�z5���I��#�q����9�j�]��O-i_Q?_�5��F��`��阽3"���~c�j�QNM'e�zc��'�)R�d	�v!��&I���UאS:�r�Nt{%kx��|`�t2��v�E�:�T��a������j���c���~l�Ahzʶ/נ��	������Y��a�!��������ҥ�����C�rGA= ��4'ۧG%O�����:{�_��Y��k��ZB>|Fr���}rAx�����H���orf1�t�5��y��;�I��iE���z͵0�|��D�{`����7�� 8�H�\~�ʼ��eԒ���Kv1�Z���3�BUɵm����wNTH��� U6;ܛh�̫�F�k�j"�U�O�'7�@�~i�Q��_
C5P��g�N��܈��*n.+
W�5e��bs?�E�}܃PD�//����������&~���Ge���A���W��'5?e��&��Kp|?�Q���<��5z��R|��c�֯Jϸ�������M�(�1��<�3�^�ޡ�6����
�m-�}8|��U9r4ʑ�|bà���B��Nf��W���dh*�Qn=��4�[z�9���b}��%�� Hg���L��;�f&�Y'*��p�ą�7$M� (��g�53ޔO	U�)7_H�	"@ӲލW�^�mko���bYK M)e֣�V����D:XEYm��^�	>�M\v���qkE��2���1�r�R�H�%��C���s.2�<����L 	�����V jv\n \_�%���0aeO>w�.�CdJ8gr�S�)���U��|�M�&¯,/������@�+�5�<�W�>�~��iG�����B��{R�������4�{���7���JB�m��#+��}���D��..�}?���b�Ҳ�}��)}9W;�iR��4n'�hH����?^��^l̃2�$r���`��r�Ht�b%_�W#�	VlWA8��F����J7�h0v��֨����)q$m�ھa,���������{(:�̸���p�Rlĝdy�1b����݁u
F�!^��-��6^�
�OX2[�V���p�� @s���L�E
�]����{����z����u�ҷ@��L��*�[~T~�_��v �*�D@�|��UѲێ���ս˲���S����o.��c!�3����y�@�/v.��F�u�۝�
	�SS�ԯ�J�;�&,B��x��k�Ryհꁲ��*�h��%����_ō��or�3����鈪>��d��J~�~���C65!�(�
�g�[!4���<�B��퓳���`��!o��C��'�X�@���P��1)�9�H������6�^i���-EQp^��C��������3�m7�7���I\kF�Y�v����
#]%_�j��A��8g�D+��gޥ���D�/=ԙ,�!aml��% �U?��7��q��r^�Ȑ��R1�H%u�E~�@Dݑ���l�.�Y��_,ϙQa�(kTa����<����R��#ۗ+���}���ܧ\3+��ӷ�ZA�����Ӓ'�<��
~���YlQ�|EjF�-vĀ���q� ���}��^�$�;����UeB�#�r�)����� ��N����Ln��]ZF_��2(��(���8M�mL墰�㒟
)y�YJF�hN]����	���<�U���@wh�@^�|Ȥ�����4�>pSEv�Z�D�Y���_�T�v�\��Ѓ���O�ʩdUS!^<7�-�$����Gs���/��p{��R�,�<��,tt��<�yx�X�U�tS[e9z�Ǭw�5�J���gK��z�ʻQ�
w%�0Σ-�ZƼ'����"����G �9����v�b�jl�~2����������왻���t2ly��3CVF�[�*�W��<3�/fk�К����)�!����	�`�̈́Ɂ�bӫ��٣S�B��2j�sn�E��)^i�#��)Ҩ�Qt&��OL'ʓ9�W���T
V ��!���zT&?��(�<:�"�o!vv<�����N�gٌ�f'x���s
$֟��/�t*p�	m��d��nH7<I�y��j�O^q�XCi�3F���\i>%�A:�]�Д��嶥TJd�?-O��}#[�x��C@Xύ��lg_mƑ�!�TP̠��ْ�c�o�{�u~�H���x������	$��!E���P��ؽGDU��ls��ܷ��G�5tl�?��o��~�*�X$�<��ɉd7;��"?*���>���e��T�י{��8�w�e�b��_'��%ÓX"a�d�M����a͙�G2Yt7���I���UG~�gÊx�Q���B�0ZX W0X�$qT���8�X Z�=��j�Y� � �
� ��j��k��֋�l��s�j�㨞�k��q5U�+�;�c3Xݬ�� ���#��t���g�v��T-�?k�q >�Ʋ|g�@�
����
L���xy��%ǘ�'�L���#lFBO�͚k�mL\k�)WF�z�V�rN3��n�ֳ2�p��;t���n$ Ge2M+��r�&�J�*��v_YN��~E�q�5QلHmJ��uL���g�oJ>��@Ȋb^ƶ���-H�#~(�qK#撒��$���V^ڃ��Dɿ\Tfe�Ъ����"BEQ�a�a�ᘿ���������8uksE�k�~�`$7z��L*��Ѥ�����uL�.��ҚR�������iPj�Th��7�����\c��I`�SPk=��$s��86��k/��Om�������Q�I�)���)�4��+I�v4>�ȓt'������������1��Q�p]=F�V�/4�ޘ�[�u/���c��>._A9�S�h;�	!{B���T���(��E���YYu)SW�u9J����:�S�$Θ�,������G�����4�s`��)'je���e!��L������P�K#Pө������M�AO��i��A�����E�JC��+n�9ŪNX��1{k����%����ڬ}ì��.$�$���^|�����AK$�,] ��ܺ���@�����a��[��+�#.R���U�iNkD~�>��ǧ5PXeg��r��$���v��渴��4�Zv^(j�U_l�s�s*����y<�� � �S~+ze~%B�(�K�~M�v#o��7����
DM���:�"����W�r$q���t/I1̒(���b�lp�����P,� W��&�O?3㑦|(�c�;�{�Uc�Fl��)+��t\::9Q���v��F��j�`O��h)vIg�q�zlW���_{������Y�4W�>��1h7��X���R��&�\��Kd,'�L�g�=L�����K�mw�J�Dc� �7|��D��[�s�oǌ��������#�`����®!�S�'3�,F�r��Q&���w([�$���u�aE|a��d�P��6<�Y�8h!�-�f�]�ҷ*��t�����0~�P�kN�dK��:	.�@�w��Q�q��m\#e"�����KO����[ҥG�J8������;-m��F�'��pa>_~⊨͝�;9։��yW�!�b�q�.�,��s
z�]�}>;�� �db%g?2��@-�A�?ԧ"@`c�N�r��^�R�8�_!��� ��n%j�r���Yc�3��ط�j��0J���{�u�#5q� & �8�+�@��oATt�N�I[�(��n���h�"���y+��p�0�������JJ	㯁;����/2}u
��6[|CI���eQ��H_�HV�o���w�Grs�_+�����#�"8�98���tc��,���,�[�#��#{>��� ��%({���^t99��A�gA%V�IE�ܼ�z����z�"@��?+�S���}a5	�Y	Gc%��J���f��9/�*+����"�9�xs�1�7S���x}(�I�쯑fF�G[WMն.Uۗ�eo�<�&w<d��!�Xuu�o��|@a㫴�.��]a��XgM|�����q��Ԍe��&ۉ,�s���tBx�գ��mR��+�T��(��x��L��?P��-=k�_c���ܬ�Z���n\�3⩏�$�w��p���:ƹ|�H.)A���������-.�h�M�=P��ؔY�X��3���S�\�όz|�A;Y��v�2h�#7Y0@]{R�0� �/&��Ϝ�`�W(�T{�03d�7��B���݇e��>B�;�b�.D2������n�R�InV�sZ�ٝꦮg�r� !ZK�R��G�8a�_].�5�����Ȱ��k/�yl��.X�` ��л��u��n�s����\Pw��[���L5������Wꦎ-�j�-������(�юrM��*9��~�<V*GV�Ƞռ ѧ	�ux�����L|���`��^ܞ�8�n`ݰ��p�-��\:���>*�Ϗ��@@�R��Z�P]3IC�{�!�)s8�8�!B���A��1����!!M�Lw^'(���`��u(���Q�l��)�~~-�8%��d�X7�O�05s�*���
��Ǵ��ûh:f`��7(D q��:���b���HQ��$q�˂��M�V�'1>2�ܒ�tf\a���\v�)��Vt܊��ZYqh ,��g����>�8�F�[U-��
���N[���T@۞�3g���q�W�i&�ǔ,�[��������$@)�V�h����'��F@o���R@`tf�Јu�38��߂�ܜ4n?^���� �:�g��n�l`o�p�������8W�Aԕ�C���~�AZ�v� �gu�6�3t�s��(��٘�Aϐ��Vwz�� |�\�v�F�W�ڸ��{����W�%�{HN[�����}6�z]8��_���j����90k���Js���ݳa�[$e0��Ŕ �|��M�)ٌ�MmK%rxP�B�-y��\J-N,H�[�T���I��*��m�"�ݽS�*�F$�@�fW����2|5f^0S�f�n�-�q�a�t����*%>�W���ٱϺo<�@沢d�M����U�����,$w�$pD�Q�yB��i�!(@��<_�'��q��h�&�{&e���$�.f��x��ش���n�V���~�.r��֤0����ݛ ��V��J��l7hz����}㫤��|��Evڨ?��JvP�d��%����b���½޲�Nj`�p��f�/5%����d�w��0��5��ePϠ��C���n"	[�@-m�t�w�2wz�w4ڷTk��<�Ė���$*�'ɝ8��2k$��>�f���Q�dh�X�2�L���fC����CЄ9���̡������a7��v�e<���F���sw���@8$݌qY�O�S�\w�`˗¼���R�}�N:qh��^K�0T�2,���J�B=���'������W��cT_P fG�E=Y���*H��A�p���smEo+�hb2"	�����������}L2mrJ�?' ��B�,x��*`ޏ��0�L�t���h�L����x+.�<�OP�ٖ�<B��s8��A� �J�2x�OƳ���:Ss��d"˔�#3�$rb���Q'Iż�BWRɶi�/7_l��za5`�#�+�蔾�����?��d�;�^]�OX���֍�m��s� �����S֔�5Toǔ����x'�+P��l{,�i'�)��9le���[#voU`5��Ԁ*���B��+��	��nrZRa��"'����ڢ�N�/��5�hma^[�P�^з����6ߞ7����H�;���q^lehI�I��՘�Ä��(|���h��P ��$L�By!]w(&�<�q[9h���{��;`��h ����t}0����"jA����C�|K3���������?��y���q�Y��a�����Rn-���]��[���|�Of�-W���̗������g~%^�(���f�=��rb���5C��v��{�Y_D���w／t�����W����ſc��D�RzV�!�7.@ �:�S%�;A�����25���B����A�Q�O��f�ghk�Qsx�P(�z��*԰�"񣿡�̗�����{e:"q����"Y��h)�%3_����.�Y�.�g�����ۂ>�����ۣ���x����B):5���6߱�#cHC�pA\\w+�\z�?�y��_z4��,j��W9T"���*rw ��"]��P:%�����g!	M$3�o-��S)��	�ѝ�%�G�PY��0(�������t��H�|d����ٗ#PR��E�ۢ.�u<GteXf�±S(w�5�x�@��?�]�o�,r�݅�J�������>�`vFBL���l���GAE#©��z�o��o��I��c�9�W��Eb�%���o��ꖋ�����G�`��5hT ���+���1"g9_c�*~�4�� 6I��G3���|(�{�� `o����1�צ"SwIPx���ibd�J���	6�V�'�LIq���Qm�v��������LR�	8š�.EK���h�
w;�-�_S˽D�c��$�����߾]�F����bAr�=�>��*�i�'�#���T��c/2xi��Bшv��|l��>i���woRx�\VD���E��[�����	�Z��kǅ��q�ĴL��lm�%�'��8����uB2�B��v�~�(^+���z�!'�탆�ߕ������_r�jhU*�R(�X��;�7��NA#s��&�ⳒM�q�Pl�\[�R���;ܱ��չ�N�n��r{y�օn�_5�����v;�P~Tځ��|G*�/tӄR+8�+>�:�W:	.��<��)��~�Gw����|Mo>��Ȼ��4�n��3f
j�6�'�����D��[���`�g�5$�Њ��N�@^��[4�7�f�t`�?Mú�`_�Zb�*`����|�TJ�ӯ�w��c F�xmQA���g�8�6��4�>xů<md5|D��$���������B-�R]��}��g�[Qu��\I���~w��H�MA�O�~U�$=21��Za�&�5@=4���moh�%."1~(��h�~�Q��N�����C�Z5�Ł�C��je��dݔsN_i��sj�R8��4мF��JӺ_݋�f�������%[i�ǅI���X�L?��N������T5V��Y��O�ϣ[���E��XI�Z]����|ᦺ~`���������gvG{�EzkSO�Ж� ����5@���AoH�zE����$���2��yͽ�[�//D�ؒ��|��y���&�ʧh��4��3�Y5lyԘ[(<�"^te<�,��\?�f�d�S�dd�՛���y�'��;@����o��Lw~L��#�β����E־ʈ9��)�Lt��NH�9h�m�hZ��FO��@ݤ��9�?'����Z��۴mYHA��&T7����$E�\7\\4�a��E��p?����S�sG�$a�K�T83�Ul	D�!��=ngƞ�I^3������ J�/�Jdx�L���ԣf�nR�xS8C���Jl��w#u�H�D�J���9�)����&�a�.b�>�Rm��y5�q�̆�aQ"k�8��V탉ʗ[�"gw,r���&�_��P��.e�@	��LD��.�.<�R
�0�O���c���F�S~[i��(���|?�;D��1��u�r���a�UKF+s }��4��4gū�8Ҟ�J|{Lhǯ_𢛻m���'��!�w�G����Z*�ʘ}dG�vTo�lޟ�FKL���I���,	z� �� ��KC�����X�����̘,��اb�~����K�V�a8��"�6�[�J��W����=~>���Jά��w>���T����fFBW�Xj�"���p]H�઄�eB�aS��,'	�G��5�Y��$8t�k��ka��K%´n=�Փ���w���HHQ��m�<���"�ol��Fa�z���>|h�%�se L�?���X�m��ȃN�q�6�0DO_	;(]�K�kbF`��R�q[��ܘD��D�$%W�)�e�ZF��G��[�+(�6M��54(Y�I�v�w�ѫ�����s����x��(��(<�����>L���b-m�_b|<�j��Mf��"�tbo�{8��X��/]�G*ySʽ�!�i�5b�W�}(7t	Ђ���� ��T�@���vR.��D9�ⲫЦmK�dgt��*M��)����)���}��A��}:U-�	PW6��E��o�B���������M(�iQ���3>#�dFᛒ����\�hw����A�j�C���ux$�(�}�L9�saVL]����DE��2�aa��3���Fo��/�"c:I���N�F��A��<�(+@Ⱦ}��^�\Y^덏�	7�{�Sۧo��6\Oc<S�A$X��R���v���r�2>VL�0��
[g�R��<Wc� g��-�s\ߜAM�����
����T|\|5B ����-4P�����͌��t��v���pb�f���Z��*��u�A�c�:Bd�j�*��L����f�7fv�i��g�^��(>:l����\hƬ��q�R�"�M���3Ԣ��I�Gߑ\�9�Ϥ�t߷�Øxu���(�j�;.b�L%R.U �lTf�S�F���iU%�ڵ��;��,p9U^��?�D�[�l�}�JJ}���X�,3`I����J����u~�tL[���ЀG9��F����'B�V�mhx'lB؍�x���ĳ4~Jk�DD��5�$���"��<\���ЫKu�t��&��+�D*��@� i��DߑdIi��w�NX)X2&g-wgT,W�g#�2�� +�x9Kaal>�)��	mP-^HF��Ɖr^W���+�o�<Z�L�c�&�B�|i����`�3���PՖ5����t�ԗB�U�7~�#��6,�6��u�4v5�Xݩ"?�����a\�8��^D�G��v�Y�>�0��8N9�4�P�m�y�+�9-Hz���r���z������Ѫ����:���LhsE^�� �	Xy�*����È���'Fl���A�ٛ��x6�%�.˪~�1/��}�h�J�{���o�\m���psOK:H���cQ��C�%��H�B�i�=�@�>C��`1���,��wd��=�G	���ܟe�.<a+��9�Qs�Wy�%˨��\�����{����Yx�{�c�_&�)�	�α�Z[l6)����TZ]e��{�d��#�Et�������1��>��T�HhW�?�]���&���W����"�|��n��F|�RV�TU��Y�W�3�|��䧺���Y0Z�Z"r@-��Biz�nfrJ���E���]�R����j��h[��y�m���8B�����g���#�1ЂwD� ��/���{\�k���J8օ�� ޡt��3X�
)}ф�r��H}h�W�O<��_̳���K���/���S5v'm��_�UwRq��葞���k��տ��~�z�	�9��C�M2���U��æ�[0f[�ݶm��b&�P��i2��F�Ɇ��tlwM�w�%�& ���C	�1v�s�H%=Ep��=@������Kr���{r<*ED��)�l
2]��+��r�{$�#�R5XJڰ��'�J���9~�X�"X�;#�����$s��I���L��L��;$����OD����vx,$�)�^bk���qE�|Mi��Ӏ���n��5huq��5�PS�䫩��a��%
D��Kय��L�5�!ay����6�p��
�i�}"�K��%�x�B�:2����~Il�@ec�z90�;����@|�>-��3PdS����S������uZvXK�&�����g��L �J�ɤS����e�_�( c�������o�f���`l��5���G=���}�t�ɬ-*�{@�.��+ �j8�I6p5���G)���Y��n���Q�j֧N��nH�	Ii;��;Q^l>~�J:"����*`��`���ysP��e�͚���ӗ��o���1 %^o�`��F,�7ᄈ�0_�L��)� :1���A�ڳ2� ��ۼ�Q�����/�R:��0qv$%��������!��I���y��c~ұ�Ƞ�&a*ܯk���7�4ŞX��?Y�d�R�
���[�������u�����jA`������Ʈvv�M����b�tXə��vqǁ�����,���4y��k���z���� ;/4��rΙ���>]P�.�=s�q'�␐��:�wDz9c� j��[�m%�Q/��yvZ��(�>�;/gI�y��%`xa:@{>�m���%<`ۺ⋪���ު�N�2�r��
�c���V��.W�Yl��'O����bڧ�N��2A��\b����Ё�&%�_�$�r�_)�4�C<��S9<�����5����qq[��F���W ȫ�}?��酠���z��|�2'����/�i��eOx�r1��L*m��h���'�C�S�WF�Ǭ�쨩8lXkd��dF�x������KZ'+�-&��&5֗a�D�&[��9pS�q��J5X}����A��J�������"f�7rd�¦��n�O�~�.�hs�~0]�^�O��c:O�PvK�,)�
�b�5�x�n뻀���G!a�ܫ�w�j� �dK�;�ڋ���N0�t�ب�!�[S�r�GW�o'������MmG}A �ڬ�no��ENX���� ���?�!:��-6����%������.��3���U��P�����d�p�vs���0�����R��z2�L�?��3�0�K��n7��S��q��9Ew�����4������}t�*��y������������ ��h�g�ˡq�k��[�{b�E��|�.�
;Y�����!ϲ��ԕ=���˯d���`���^���W�Hf�F��k�"/k&23����3A���;�8�����ǃ���nli;�����>>�8B$� $�ͦ�w�9:FW�������X�a�}��
֦�0L-�ߑ����s�X�à��й(����P��RdL� ���[@}%����4&�W"ٝ �Gg�]�6�`����2{n��!�
��˱�at���&>��N��ܤbh��|>���XOֿ�P��@�K����V�Oޕ|�7�IB�a��7��l_�e��M�$P��`���w\�X�t�+]���=�$����A8[�[-Ñ��ӵ(D�0S�`��b�s�80�1%~ӷZJ�0<�C�l�wW8 �4�t�e<�t2ޚ?��~R8B����K��� ��	>+I���8g�1e��9u��3�`'��-�� ��8z�e������8~>(�6d���F�P��ga_�C4�����1�S���2�p+��dZr"y�Sơ�JХF��~����c>��]n��'y��I.��#B�[,�^���Y'&׉r�g,t!�AB��1��ԮTb��������Z���T�lv�f���pS���z�.���X^ %}v�S�N�CT����¶��|륓|�a
�[_.�ي��Ѹč+�,'��%�	s�>2���1�7��<[و۶8�����dh� ��G��Oj��[��F����jI�址�@v������'@$���k�X 7���D� J�#͈�P@//3��믗�4rK�J��]�^Ca���"e����6�~_.r��87L20�RKG�5�8)#`BCf%b��L��k�@(�,C$$j�K����ܼ�].3־t�cd���k{}�>�5��QPϐJ���L�݄��;1|y��)є��V
�,q�ǺE�.O��v����������������𕶐Ǔ
�H�缺%��L1�gE���]�%N�ʅZ?II�	�D�ߴ;����j��*�HHo��b9*j�ʁm5@������!��{��X'����A�0�m�5ڼ�� ¾/mR�|�e  �g(������W
b��"}���i����������B�#�	��bц�����̚�`�Aw�#C���tk���]�O�~-h!"�E�8p����˞�tˍl��x'�Xƍ���p��a|��r��N�͎TD)�ﶨ��tU���׳"�Hh?B~���n����l��2���ʪ�o[��_��������y�n;���x#�ۚ��ͯ#�('؉��DwR��.#T�Z���g��n�����(|�A?��^J�H�%�^�v*�iq�>���'EVS�I���~��\o�O)'���>� إ_<0j(vv.�8*ȇ��$	�R~W�X�1���Q��Th�>g/�u_��KL�<�����QI|��Rx9Q=_���@#�=Uq?/.�
�fw%U~�j�,���:!1㨘:��C��Fvhu��֜:�
�+q�6�v�����hǕ�q��E'8R��c>�$���Y$����s��`�;���������;�I����.����'�enCmpU�.3h*�(��hz$Y��ƠEH��zD�י���`ҏ\�1x��A]3�ܤ�� �k,��<L�����h&���k@ۓ�2��ll[!����A��"D(�Ӂ{i��Q�!�&撚>5K��S�sGS[OMY�P�eN�d����3�����ǝo��ݬ����s�O�˱����kH]ΨE�ˉ_��w��KEI��=�f��ͳ�5Ůfps�_��ȱ��}f������V��J���f
 /R��w���T�Ј	)��V�|;�@%�s�5]m�'B:`�l��MjZ͐��x�X7��'qU(��y0;J�fW�����k�o;�3�~���!�7�ц��m�K�}�`�-�UD���ݱ��x.�� ��iVu���n2B�,�eOQQ��s���*cm1�8h��X#"���$6Y.�ςK�xV���Q� �MGҘ�Ib�k骬��/�@s��z�ޖ��+��������lg���lC���}����b>��DC8g^R���U� �J"&���Jgݔ=���⸉�	�g�T�_�\�	Z�cAѕT؂�7���l����J;"�F\ c��"�� m+�S��1f����1�*wʈ�䇮y�����-��d:+���f#Y�O�<+GA�~���|�.ۦē�~�<!�}�����H�쨴чe���ji�����tE.�uO�F��l��~����夸�u�B���!��u�jm�)�6��R_ߏ�(_͛�O�ɨ!���d��'1�2a��[�C��Ւ��	���nF���Fx�W�4-c����<��Z�Լ ��}?�(1W)a1L٨�M$	@TȥF��d��D��]a���x\U�]i���hE\)�\^��Z�89D�+#�
P�ȃN�������#$�&Y��Z�~����_t`���5A�غQ��GD�	��.�l�0�=��PV��C�q{�� �?�$<�5[^��۷(���ɴz'���e�o��3hʩ՛��_x�[\�bؗ��(s��4�%�t ���?�kRS�0����*��))X�Cf��7GtR����߽�s�ܒ��CƊ7Riw�/�$.���D�O���|��SeU�\���o�^�R� �,���<�������nބ��&J��ޠ�U��KP4�J"N�*����ewK.�|/���:M�V��p�yz��7�䛴6Ss�<�^���:ot��-�G��x{���DG"q+��ړp��*��Z"��0z�f(� ��#	M��-�'�2�iu[V�[lAg���@�ayv���`��:��@6��]�z�}�BƳ`k#v�.��ā�̢�w��$��W��L��9��1�����ъ�8�~%��I�4kV���"pR_��l:wd$a5!��Q"��ةA��&7�΀��VX�����ۯj��!4:���X��9�����=���P��������K�y���L��7K��i�<#�J�9Icj�2%c6�ۙn>Ղ>��excRR������qMd�E��vqŵ�^�¡$�R	���|j��)
����u���ˢh�a�́W1�`]�L�HiE�q�$���4E��)�5�J�6�ô�Z+fg7�T����O�jq'�>/3�fӅ(�i-Ψ�K�U��{���rY��=��W���6;�:>��'�`ڴ_#�_���K�	��e��Cal՗��[Fb�W�%��2�/�|z��w��$ԯ���, Ĕ3e�8��j��~��ش��xY+�����b�
e����z�^�^}�S���M�������iK��Re`bǋ��h%��]y�%�'�~�"���|�c�p����Idzh��Q��ͣ.�rX�`፠�e��#9�Zfrf��-�����?�q�pμ���>��k���X[m1��4�1Ҿ�8 ҝ:7��~����K��(��0qc���3!0�a�LYx:��y���[��}̈́u;@YI���.χBX��e�2���h���$�5'tj�iv���x�F@�R>ͦf!�ib�^d��+�='D����P�,䥕<yRI��>�I��?q�fo��;9J!�����Onx���ad٪�l#E�;��"EW����!����.��c�HT|Z�r̡�5%_�뤐�>$3וpe����^�/���1S�T���Y(#�v}����Ro8�B2jy�"���.���Ƴ}�k�R�-O:&��n�	W�}��6Z�@�e2���}��gB³��7`����V�Enb���&įߐC�F��Mm'��(S w� �����3�,S�m����D�:�Peӌ�@�ޔ���4*�%�	�!���~�3!Y�C����K�C��ї�9O~��a��qK'2��A=�{#�HD�q��I~���Jd�(f7�)��`o�h����Vg�I%#�� !�h��K4~M!���ȕp�3�I"�Z֏����)d��j�){'������b����XX���qī����˴nR�<�H�y_���vR�Xr�Հ�qуAJbH_%V��}>�4�%&�x�{<"�mh,�o_���k/�*�����p�l'�vg�	�}�p���S���}AUL�j�:���ck����n殺!菱٭A֪�F�g��?��5[�*OIg~Oij���%��4�'�usxj���#K�Z%��}n����46�~��+^�ӻ_��ǩ��W� �ܱ����{�ajF�$��ы="��iL�x����(���)�0q���=1on���̧;��	��G^U��5��^�n,�K0-L����7H�"ݢj>�"1C�Bokq3&}��a>����.U�Iڝ�j]A��@����)����פ�?��$b��e˞!y��[��#մ�fܓah(j��-����D,���7������k�d���|�w����)��o㰍�Q���&�a[ m9i�(�BiI�� ���h�7U�
���z�^�-G�_��?��Ju����fgSN��^�r 3��
%���di����zd*?���DB����#S�����'� �B!���H���K�bk)�h|�Y�Ѯ�X�6�c�.0���H\@��*�N�0��Kle���u�%���v�Bq֬9��;�
"����F�^&�v�-��?�I�$���k��lE��r��ぺ��G�$&G�{�2�x �aM�#�v�RV��[&�����V�	�����ºyVr�N�o��>5(g��BxA  �[mc����	S���53�$�u/b{Ty�m���6�c.����_����q_15�B��u
���}���� N���ī�ӿ������~B��9T�K�sgի��"%�����Pw� ��o�O#����\Aa�9H�u-�G�5��Ƌ�����NfW�C?)J�C\cW ?x��T�>�+V��k�|�>�3iS���ٴ�LeRڔ+պC���Z��9�Q��tc�6�DGNM߬�,ba�7a��/�l(�D�uL�Z.>wpx����R�0P��<F�i��7��n.m�$��F��)Kɏ^�rΆn���j]b0��w��yLr6���h�OF�?��	��h��|F*�v��Qc|w�y�"��EI�90�;���D흲[���Ev��.ȿ��"���ҽ��N���G�fD��ik��D|[s�є��.=�~10��,h����	�rȯiĞ!��9����]�O���>�<OtG�г7YW{GN&�~%=lO��A��w����JU�Y����$���*���oś�h�"�d?�L��6}�w����T�˱`WD�Ѡ���ћKÞEI,�R��?�Q�Q�A��������p�Fx�x��������A[en���-�E�xԧ%�}K��b���o,���h*Ʌ{y�)ɫ�U�#�SH�j2�����U�W��L8X���n������p�jBp�g7�#ް�7�	�}y>(-�~�t�3�RU�WF10,ǳ���S�X�>Z�_��_��5m�|��cD���H�[T�Y�Ђ��d�-�y�<Ozn�~ ]X6��$�.G�c�fzM�E�d/�	2	/�̨�o�L�Ͽ\ۃ�m�Sx��I���+�f�ɐ础�I�%@gL�u�{��u�i���OR�D h�w˸��2d�-��-.l���1��(
�����ɸ��O�q�n|�!S�7��	�I�ťG�!=�u̧�����09qة�6�����}#�Ζ��C���/庥�z5�.�\���U=3ge1�ac:^��,�}����;�C��k�.}�|09B�+�@�v.}Ӡ�pu~�B����i���OH,k�B�.���ĳ�W����|�G70�|'w��Tu��.������b�w�0r�R���Dx���kV`"�`VW�fOy񅪘�pC�T��Y;�]66���-oH��Ǘ�Y!���Kz�u��=E�A��"��ʳdl-�1%����\���f�X�r�=�e�Hp����U�k�9[�`�F!�V�k�E��2IO	�rq��(��b��Q����\���-v��N�V����l�T�'[�BZPa8Q� ����5�&S���o�Xg}pj��;��P��ɿR��#�O�X(JSZ�@s�����p�a1����d��o��l:���	#���+�� �ͽ��-��~L��c^E~� օ\��O �&��������E������̹���ӻ\j�"��3�4�MS�ָb�L(|ŬW��Er�	����������p61og٧����/xB|�n�0b���:Zl��ż���%�U33�:&KЦ���iuʧ����?B�W���hi�&�|П���3`^������76>/�K�\�͞B���HTItf���|ᚿp +K^
qzIБ-ܯ��]���W�]Ұ>�B���t�bd0}_,���u��A����6(8*rx��r�9����5��%.,�y��PvC�(rgQ�?�O�'i�3_7|���Ԙ��n+�%4�5�M��ՏW_���mx+����/xG9T��#�(�Kw��s?�K�r��b�ߍ��ʏ��ќ�"�{D%Xm���i<"*K�o%�R��^l��ae��
h�FW�7H5���}"ԏի�1_x�� ���E�_�;������Pl��;	��HY��*�R��?�\�0�B
F����$�Ob�#7�}KF��S��V�Ҁׯ����ݽb��h�5Jb�17��o���7g���,�ۗV1�]��ݚԨ�T��s�	t��������H �(�<���E�Y���0����#ח�D�� qV��DR{׫�:��G&�^��	 U
��Idb�V���b
�O����o��:�,Hܵ�3�4���~���0PB}��R��%@����_m�m�)�Ǘ�}��,વ��z	�h��
�S���#��|F�8�-���U�F���ȏS`�'��o.H�f`�Lb�h�E�A~,(�JWJ9��ʺ�IL�X93SqZ=3��4 ���V$B��IK�a�GP���$^n\�]жX$�bŞ|�*3!شO�<�6ֺ�CQ���X*C:x��u|��i��|�`��_�∇�$&���J����.�=W��!��K�������	k~�ߵMS2���������
�[-�k���'���L�� ��si�*���:d�IT��P�?f. ��#P�����e�̪/�*ߊ7rpBe�3H.�}�;i	�0��"����dU#`�k��/� �dZ����X��m��~.7=Q�a�����/�Z��`h��?(�<XM�QM����ET���^%ޣ����������7"��sq-��SJ9�]�~ӻ������x�����O�c,�y�+d��Cq�V�Lp�O%:;��1Ͻ;~y*q�h�� ���U\VP��e澮�{K���RJ��?2/�❤����u������DO9�hb�������*��b�rR���ČL���޺�\�@�.�
TVX��
Ë���m�3�����|�N��!kK0�`��X����q{�4Zi^[}�R���\�Z�ߔ��<�����7}�"I��|���_ݬ�; �rM��>D�ؓ�L�� _=��'�5�y��ž���.1S���	,�B�6�[�<�%�0BD�F	-�Gd���d��U&'����A6��Y�*�31�z'';�c��,aľ!�x`���}/�����[L��t�Ju�������j�R(��q�K$�~Di9���M=3]Uz���Z8[@ H=ܹ��I�}0�zZ�4��_�<�1�oxEA�@���	��<�PJ���r���jY}�Ő�w�翨G~�u �;"5�^�c=99v�⮯�H�HB���B��u9�!	�~��z_ځ�.]�0�dv�2�X"4~5���H �},y9.�#��pw�f%�
�L��}p�����&nJ�2�hR�xU×��"��������XᾷW�;�]���#�T�^� ���V �<����L�����nsp��W*��F��!K�-M��3=��D�Y�Pn�*v6nU�ǉ%���cl�
̳��)d�P�@�j�D���w�_�>jg���&nu�ѹ���x�:r�
P����Ԟ�V�)ߑ����D��Cej����$�K�ܔ��΁���z���&áѺ�����Y����P�0@r�&� y	�lP!���or��xk�Oh�ØB�����6�f��F��_�It��#螓:�ho(��3����_�e���s����P�!�����ǡ����6��p���m��j��q����3�YL�����8<o����Ƞ˧
�ł�;���>�<)D턭�cv�s�?�7m��@���,��1�ŕv��maWIr�.�Z��� ���͆,
�&FF��Qf�"���)5�_�6�Kb�]���Ub�r3@�ܩ�������8i����R�\\�~&d����oފU!iP5����Hp�	Z�ѡ\��&`Ԃ5�o^��������@z���}%�J���@Ndh�_,�/�c�kV*\�z������4��:t�`��X���,lҠ�����Ӟ��; +o+���+��P� 1
2';�~��V�B��gk�^��� �fP`��B,��52�?��APા���6N�l����X���4���#Yz�NΕ�NX�3�/�T�^�����@
���i�/9J�tY5�P)��Wx*K�^���Qf��������CK�U�p)��W.�F�&K�5�e�V��1`/u}��2n��t�Kc���5r�U����4�.t�3e����y���~=z��ON#��Q�m��%�bt%���j�EA��9J=ڲ��/P���1�C�4l��Kh�r4j�$�߅�-MU)�.�o�>V �톿GQcoǙNf�e"<�3�:�M�~�`}��<��s���W��ma���)t��/>�|?�1=�Q�ս2P��<7,����b	�t�qձѠc��bõz�����rӇv�e�w	]k�5� �V-���F��(j;6a�%?���X0��H�Z���/�:�k�)ɰ����g�m����	k>�u�x^!�񍦆������s3$Q��>J{��6p% "��R����a���{�vL^8�k���0�x��P�юL��?#�r�Q��&a7w�$����Pjv�Ѯ@�q���[�bb- �����aeڝ��0,E�����M'3�Y�I�̕	H5�@v~յ �<�+�&�0q�t)LN���Q�x��QЅh��d��%��	^\�V&�ͧ��m�k�L�_����5�v*�����:�_��"EԢ���smk��$�,h? �Ϯ���WaN]��rc�`��(D`.s,J�?Bc�!F�^�6@�s"E�7�f�������8��Gc�6������E��a^>�a�����*�A3���#Ѧ�`�}���n�ѐ�2/��&�V�e���.��weU���xƪ�s�ޤ ��*�rR�K���r�WQtV^v=d�ϟz�� �O�+Ѷp]��o�q�{��1?��uߙyjr:�<����8�;�������ܚ��g}x�[��t���ј͉S��lKe0]�EV9+��*S�cX$�;s����_��4�d����+<7�� �R(�J1O��\:MB��6;ږ�9\���]��Em�?5�aKwT�?7�����m��J1X����v�d�/�� x���v_��G����.�qcY!@��&12�*`� �?@��<�:3���wN$8�^л1���Uι,B<�����`��N���+�p̘|��{ku�焿���Dշ�F��^.Db�GM�T_����$�B�·��Nv�;��'R�Z���;?�f�?�?�ed�6-=@���`�rK�U��f��+�Ҕ ���I3�	S�B9�4Ǵ��ƍ���MԪ�^��Ck��h��F��Ў�Ȫx����ȍNo��b�hE@��AfΣ#�T�7���}#{QM�X�țC�����t-��#�Dɸ6���V|&Ӏ=`��^�:�%[����f~�-�=�����O�h>�eX��5�˫�����5��5ҁ��N���P�n檄$ ��R��>y��z�怀�؅�Tv��KR�n���<Q�c�h��@��T94h(���$�I�c�a��<կ(V�@n�6m��`"j�0Aa���s�����݂P��?ɚ?�� O����R�Tn٩��7�j��o�Y�5 *�iy�@���w)J2O��9�==���:=)�m�]AM��.b�B�4 uVxs�q-DF�H�����}�
ٜ"�bLY@�B���ڤ�ޣuw��h>d!�X1�V��Z��c��I�U�07���/ުW[L�/X㦰\�r�#8ٗD���@w�a�q��u=�E��P�6�NؖČ�>7G� �,x~�	��(ԹH����Jap�<G��|g��'w��b7�^G�[g�t��(�?��cP}4Vy��9�*2+�p�L�J ��㊷���h��$���=wh-�~�?�|�k�{(���B���O����f@2�i&\ �x�$P��$$u֑�=lmbv�>ܙm�W�5T����å�Ih�~��UD_:�B�#��պo�$�vS{�&N (@dٿQݽ!#�Z4m�9�-����q�BJ�8n��{(�����x�L��l�e�o�X��tV�ز�Cf'���2jmDtq���,/��hT����SބP�zCߵ�t_�\�s�-���f�H=P�\�<��8���T��>E���ҧ-P��~�a�ט|�N,ڦJg�F�s��Q���j���~Ԗ/5.7w��YO2:��S��w��b8!�p��_1ܥb��Ҝ�Zy��d���4�AAQ�VXg�Z�H?X�T5N/�5�	xB!A�*�X��J�XA>>m_[��ٝ����Pg2�����[�h�F��C/LZ������~��j��M2�n�`�Z��g.֟��D�;}!ט�M��W\IF�n�a��eA ���g�Ɏ��q���m'����f)�G3s�_�X�#�{!�k(��-��F�v�
�!Ϙ��+��;,����=QSDzk���)"���R���ҍ���ޤ@�����.�=r�Uo��aXu�!�� l,Qȷ#���)Պ�\����DƁ���\-d��T���u���	 rǗԁ�}w�K|�ge�y���H$ӏQ����OhO:u��@��
�tm����#ZԔSٟ�����@M�XEv���.S(�"6=�Q�,�6�&���`�~+���t�MUL.�i��П�Vk1s�3���PP\!�}�An��Lv� P-d4�+#�f�U�������T�[����(ܨDϢ�I��Q�_$Q�#ix�E��c��;Ph����~d���#��X�q,v*��P����f5Cm`u]�h�sn��)�]v������1^l�mѷZ��������s�]eR��}Z�jx�ȍ�0j�8a3��G��&������n�i��I1�{��f�����t�\��q��`҅��[-- �7�Q�o����a�/����f�.cO)��B�W�Z���RU�����0,z6�����n�2S�%틞7)<�x�;BYn��5=�jJ
�p�χ����D������^�r����ɝS&�zD����w���=b�jͷ�KN-%0���6��3���zJ�#P� ��3Kd�AR�7�C��$V�XTt�:^��F7"���^u��f6�y����V���h��A�j���9P�1� <�6�/�F�|12;0>!^����Յ�^�K?r[��N6������ƺ�r�s�"��R��|����.��V�·��Θ��#����k��s����V�=����k+����<��RV���J\|`_`�E=]J�y�G�S	���e������Hr�x�X��C����n퇾1O���/�qG#����:��9 �u}�~>6�]~��)�ѻ|K��ޯ6-{aZ�� �yO�P��Р�|�n�{a\���	�vқz���q)�ڊ�p�L۟ٯgp=!��N�]�B�y}g.��z�"�������CZ5�~��c�@�;"h�IorhW'I~��E���~SW�� u����ʣ���aSo��LC��}�c��-1�����4(�x�|ٛx�����Fp�U+F� d¡�H�4�+�w�1eRߐ"��]zM��Pn��9=�PL�^�x4J��TN.
c�)�' r�=���A���?�����p���_2ѯ��9�d�g�i���`�"
j����tևq�!Ƨ�hV�R��(
cY(��q)�a���ܐ���pf{���Xte�9$M�|�|.)#�������i4�L�|�F5���GhyW�D'�Z
+��أdƬ�Ôl�S'��;�d>%h2�R��(�L�]c��v:b�$3w������p�� j/X�jR9�S��Q��L$�zv<'�zń�뼬ړ���!�g������6=��Uzj��8C���:)}8+V��4����4NVܵ��dÆ
#�x�U�M���ep�v<;=^�	?M�d	Q�T�Yʫ���.�11G΢�����
��6tb�'q��^����H^�
Z�g�pM�m�F3�?-�ԩ�RU�q,�٬2�-�=���UG ��hתȵ�R��'����Tm�hp}�����`���b�I����5�x�VU9=]��X��	�� +�}1,,�քA������D�"�8��A�<㚥�mG���{��8N]d�v�5(�|*����Q?28(c㠳��bO��i|�Xh�Z��؍����(fW r�q0�=�$�"3�J���t�Ì%��g5=��1��c1����Ft�'�_���a�]+�Hm���&��v�/������o��Z�}�~����l:��tULӕL�惢؅�}0w��үNv_dڸq�tj3��;{�B���-�<�C�ALʝS&s��W5y�uk�E�R��p.�5SjJ.�ɇ�8�X���H%�S��<�~Y�!�n]Е#��;.�G'�P�m*D�c�~�Ϭ����릮o�Fa��c�`Z��^}Sݪ�[6�������T�e�����	~uÐy��� ��q<� J�o���wn�dݎ/z"a�Ҿf�F�} �11�V]>(�W@O� d��3/���vtE8�G�K���3+@~�����$�J�5۟����Iun���a.Wb9Q\Rc��`�8��V�B�b˟*���>��^��eZB5)�/q�v1��>~U���e#Lc�����ҳ���@�O����aB��T��7sG�c��� �w�S�hXUL%{@?23aͳf?�-�V�Q�;N�O6���pe��+2w�8G7�hK1|�a~��.��4��t���&��UZ��*�(h?%q<�����C*�H��_1��"�t��8/WP��,���5C�rhZ�Г��U���M>�|g��3vHѰ�<��-S��"���3���<���]m������H�Ö��'�=2O׫�Q��=��0�f��w��j�dZYƮ߽�XD�@���p�@@����_
�d]&�1���w��N�`�^I8����x���v.u���M��� ��1�fk�9�H-�Nq,̋äP�������6W��R[g�c6�iFDpF;e�閲+Pm���M�:X�>�nRaX�M=�d��ӻ�g�����z�C��S�Z�fb�8K��RW�e�l�S�d��c�w�*|�h�Z**���#�2����O�럈��[�F�3�I��/v��8#��A��7�j	�M��?��e�N�<`J�V-��y�2��a���DzPt�,���p@W
a���ָs�+}�X��ݹ������n1^�[�ʒ<ם�d�ڹu � �+��ݿ ]	�w�]Ro����S�Y�̳�c��+�^+R���H4��(�l%�e�q��@�������]���H�ؼ^!?�����P��F�uN���ڡ,.�z��ZϞ�ޘ���B*%�.Ս��k�D6�y��k�l��LK�&���f
e���-g����*��y�>����f�/�� 1��C 
����d�	��+��vە��Q:�~�<Fi.��(�/*�b~>*V��e'�����y�.េI=q��f�<Hf�����Qt��_��puf��^z�G�]z�w�;1R���_��{X<)ٰHG�lb�e��ן�|H2{F��|�d��o� "��v��_m�4����Pe��b�A��{�I���̕Ѿ� �g���އ�h�omS?�hI�>j-~P�)f9�a$AH��+��Q��� v�o���UI/щ[V��!|p$7z�E�Q߬�@�Z��-��H}D��� P��3�g�G��e<0�fR���~_ם�|���a3e+X.���c L�E��d��M�qH}�-�,h��%���ѓ�#Ww�|o_g��
��D�E��mԨ��y�N����D]�Q��7�{9�´� C�u��c��>�[?�d�'���%�{��~g�V0�)��+��Oogt�)	�;-Lv,��α�ʇ���8Q���|�,�%S�JAo ��I�^�:4�
kes>%L��F������l8��폠]�/!�x� |�1�QIb���60�P���\�)��z�� ��:ĝ/M32IG�O()�d(jGk�q/p��O�t_A��h[�}�UȞY��pȋ�W/����NX͢�o��:�u�8�����y>K�6�0W~�s�{(?�.�y2)Z}	ӳ�����]�d��8��@�b3,�&�l����sA̺ �Uc��\ǐ<��S�j;܊U=�R�u��;�A��[6��i�<Z�{��%>هO��C��@*��B��5#�|t��ꜣt;`�#u�.Ž��Ř,r�3��P)���{߿A=�I?���u-l�.���;4�	��Wo0H��rePӀ�۬3�x�Q�%��*nNg)��W22��^r��1S���Y��?YÞn��bB4T0<A���T��[g�ֱ�Ӝ��p��J��EJ-��l������ځcQF��G�F�mr'�>�_$�DCe�/�� #��Nڡb�H���㹄��}F�H�Л����s�}�V�D-�0�z��C�2B×���ͧ�� �f]�y_P����F�a���t��Ȧ(58D�.w5������"�Ʉ�S���4����������4�֘/]CmxtBG∆[P�ӎt��5�D�IA��$h���9Ro�(󿭶�¥�����D��:����/h�6�Z�h
fUG(g]$.�74������Kd�,��g?�
~�l��ࠬɟKd;�oJʬI|׋#Ny�>�),=G<��z��uM0�=�]f[<��8W��*�������H�2��9��E���2BJ�|d��/��]�}p�x5l�{97�ZE�/�y��t7yI�;nO�I��#v��f�M�mJ�n�/��S�Ђ�}��ک���59�B����jy"`� ���忊e����*�'~�7A�TEX�,~�E:2�/�`�"���!��Y	y��} ^9�o��1yHϸ�ܯ��2�A*F��x?R{'~��ɖ-����=�77�gf���.�"��#���۫����z�t݃A��3"fp:�Q�_Hw�W�F��KHs��!�p��Єc�:��-ꥣ��Ɗ<*i���a�`���'\q�u� �r;�t"D�E�{�0�qY�ݢlpti�! �jcj��&E��.���ܱL�'k5L&�Y �b��\��d� ､B�St�UMT���cA9׎9�g8�}�xe`/g;#��Y@�3w�CL_u���nD�F�[l�1�Cv�H��8��y�̳y�;>��&P����%=�jT~a�U�N$����$1Z��ۀK;��o�C��y1h�g �[S�B��*alIV��]��+���ð�����'��V޳�:�u�~tI �������f���%8�gg�n�� [�Fe��"d���^����`�]�� -cR�:A����ġ�%dF����9����!�O�!͆6\�Uᬞ�+�D:��5��� ����(1Q��#U]V~�\:�@lV�|`���gC�Л4<o�ʫ/R�zò�;Y���F���qa���}��߫bġ�>�3���^(�D�1�=�'�G�q4ѶP<���N��f�	/;��uR�k'�k3�@^�d4�����v���Y��/�3G��	M'��By�Gs2�ũ;Ø4�,�D�[ǿ���$V�*��TʖL�~K�����,�I>%y@L(��]O�	aB`�6D�5$6iJ�#E�R;a�'~��Yr�6���Λ���<{�A7=Ê� ��D2͆Aa��}��v�4g�;����+�Z?m�Z���l�7�9�5�+�c95��Q�GA��p �ϖ#86K9	9[�>�&"�KU84�}\��oh���!��\�:���$�M�܃$����4��������=�W���j30d����	�S�9�C���#\ޅa+������1�cB������D���сG�G����4?�Y���� e�PU#^�T$R�D"<I\XF�'(qٗ���K��.�Fj�7������G!�}=�g��o����^���}��ua�ϓ|��(�)��׸+PCgm$�l�7w�+\�f����L#Ɵe����/���U\!��)ZoH�ۛ	�9;!��P���B�gj^σ�Ō�$GW(�2'>���d��R_�ԧ�"륟��)��#=�H;�r(�߈��;���k�|�{���X�F���7���j��х�wxXt�5�H�D,\QT���	�J��%���f�y��<�0Ǭ��HF�Ns���Khd�E���\�J���^�!���s�e띹f-^�j��^�n��'��A� af]a���-69't�+v./:QǸ2Ĭ��ڱ����)�=v%��%�ָJjg:���$�Y��	xU��K��~��F����T���؂h����Pnܿ(�'�n,���É��׵�e ��*��{�,>�tY$b�.�Bۚ� ��Hn�����s��� D�>��!�yM�q��n�9�9(`���}j5Q%�?pUW2w�
Kgy�MtB�Ykj�Y�%��tĠ(h>r(��R�z�3���FjG9����� �����:ܢ\y+#~uOSy!o��zn�dB[e�b�u�JdĲ�֝ k���\so?ʹ���mt#%d����h`L�eM��b�'��\��Lx)Q�,�����Z�_�-e/�PdM�G�m% �?C�BGC�ܷ���a��$�Nl�Y;~��ZE��4J�y*�Fn�<~s���B�����1�C�ǒ܃F��'�����oyU@n�T ��y�c`#���Am���(��٬D5S߶$��W�� �H�x��y秲2+G��H���(�MI԰��^�lT�����U�t�TOmw��v	c���lJ�K��A�.��d��>��`� &�{���D~�(���憚Q�=yn�R��vlY;�����ca��kѨ���V7��vC��)lo�G�����2�����ܴ��uK�V�|;M��/'%@����vC�y���
d��<�����ڬ�yl��L2�	�a�n i�/ 97���o0�f��O����XBb2����X˷z���	}.�)�[('+�ڙ���j�$��e���M�t&���F*rl�F*NAZE����%*�r�zj0�A���y�c+kg����ɺoA�uM,���f�p//��?Gɧ�&SH('�,u���F�K ��ZQ�V ������>�e������~B7��T��|	�'G�Q��.:I��=a�5�n��GR�{>p� 6Mn�������p��\m�D�Zo�翭����gi���QL���+��.�C6/ʮ�,�W��o�a(�t glˬ�]�n��I�%N�ҭn��BS݅~����!O�ez�U��^�}� ���6����SθϋVc_���;t��%��η36 q�bxR���ZO�<��@ਜ਼ utw�s )
�̼�A�:�pAg�������S�AāV�'s{g��j��؊J��OU�[���,�������\|��� a�E���i�.��0=>?�%<���>d���\p�0�B�/v��:߹��pY{�Rd��C:�s��)��et��F��bx��X�Cv�\��uj�h�H�Iݾ�Cu�"���^��'����R{���d�c Q�k�5JiZ���"aނ���!�H�=Y>W3��7�mzK�������U~i�H�ً��K�X��r>��"��_�$�b��WJX�Au�p�g-E(��۝����(����I?����ԫ�NvFr|�=�C��)����_����b)W?�('��7!�f�w�>��/�bb�� �E{֊�f9�G�'#G�}���vg�yb��Pq?�[�WΧ����G���#�u{��L-�*\�n�N�̖���� E��MD:���]�(��[	��^�QF�K��+���p�ry ���gm�E~��|����� ��KW�?3W��} 9P��|{4��T�MahE�n����"�uʺ̽�']�I�U���u��G����{�D���NR�J�J��H�(~�o��YS,���Kن�;I	���!g�lj��\�EW�c���¥>͌�*���+�FH�Uy���. jp�!���:;�SY�������2��|S�AA�@�eW�+]�^�J�z0$f���F�����]ԕ�.*<�mɆ{�#�e��EF���A�r�?�� v�Z�A@
��i��Z||o����g�
��y���t�X�����ǡ��4�`�y�^�B08�cO��Qވ�������H�䧫�s��������/�x�5K&�]3��w�s"�����L��Ň�z3j9j�at<<J���������e���T����`y�%w>X�6�%cYݪ�x��y)K�D�{�bU�
>�@��>�׼���G���J���֣�c$�D��ۄ"T��I��F^�p�n��D�C��S �N�$E^5.N#�R�嵇��.��E %˸J�kB̋t�Q�G^�P˳y��X�����ˮ�-��B�o��1�"����'1�� i�?�y8~0��Ԣ�;~��8��K�D��Xf-��^�s^U�ț>�v�|�"k�B��kGY��{(�ul*�>����8�[��k�G�n��*�+�����7��L7��zϙ
7ܶ$��FD���@��^)�.nsԡ/XFTZB16��h��$���(�W���E6W��\Muk����G�U�w��H�2��֒�bw�=�]"�<4���ֻ����.�J=P���y�H!�͔�W]4u��n�J�Ʋu�G����|�a�y�L�;��8����2KX!�w$�ȓ�dp;�e�����z��L��;�Zp�kvB�c*�L�iEnYoX�R혵��ܤ���xC�U�f1���0O��4MJ����"���)b���?	_��Ԇ9Q&��)�d�̶��zj���qp@ѣ'�K�����4bA��C�
[U�2ã%=8
^}���N��������W�;,���ؕ�P�7�	�@�^�S�L�\ k��r�>�5WTxb�@��b*�y��n6��M�o�]����:�H�:��k߯frB=0�a���.� Ij�������x�D��ҿ��#���u�!A(��]����*ƕ+-Ȣ$=�z�ƹOe��⫶&��p�o��A�x�5�n �c��j�7��O�̒4#���L�B��?�>ȥ�F��PJ������v��Y,��P���
��+>G�o2��4h�h�fN�톙$��(B8oќ��.�Q���Յ�&�oA)�B���`پ����� ������żʂM��?M��T�0x���R�C��;������{۔U�f�1�i+�J�d����L_�����5&?v���Kc@���(�$��sv|���+�N�v��w��_�ߜuh��N.���4R��9�%)�x	�@Th�2���U8a��Y�G%�Xր�a�B/���Ӛ~oX��MWu�-���ؤI�*��%�{+���`$��7	�����}��5�����;3^�E���(�׊J/B�h���ur�/ �}���i�f��sIWu�G�nГ��C`e���x+X|ˣ�us����o��.E&"C�����-���A����m�F��&R=fGA
$\ch��_9 ����L����>�ն�[���ߊC��MW�����=����}�B������]�,y	�b<B�u���?���6�˴{B.?f]����D���Zμ��a�I��錚W�9��O>��5,m_#��j�I��CR��>��h{�2`|W?��}ܪGH�[P�*����*��+0.���^4�C��� g��LY(T�Z�1�CT���	-1u�3�dtm��:�,��"����.	fc�S�r��,��Hb���lG�s�Z4>�J�:E��k���{��������e����\���.�&H����-�0TZ���ڗ�!�p���B���1�Zt�7��m�ó��VyS:��X����XY��R�N
�h�M�
9��cp�uf�'C��"{������y����i��*�@x4�)�V����_�D;��6T��q��s0)���8�U�DPP�j��qX,��|г��˟�580Y�'/D���O}��>�~+��WK�5����@6�H�����9����<i�r�E�ڟ�ڑ{���b�ji���;;O-&����pdZtޯ�Wxv��j�F�c+�i|Wך���gm��18�?�M��_$�l?T�U�ˏ���%b��p�8��f��0t'`�蔎%Brs��W1z�ns���dW��<���ctw'��'��"(e������I�:��)�Wo�kY����l�b�Ju��A��XN�r6l�hG�ҹ��oڳ��e}#������c�y)�+�LN@��X�3�r�3�"��o3l���U��N��vn�U���<�Ɗ���\����K��/�b/>�V�&�p��r�j�R��KJ���<�t�ZK7� ��/�l�@Ӣ<K��w4�>�S��I��WA1t��cc��%����0��g!��D�O`��Ru�������a?�xow~��B�A�6˂Ϲ_�� �cΊe\�em޺���ҩ37+�ݳ�#��;_��M���N!w�aO���O�̷(
N�x�D������(`bz�ж�_�wp$��4��#/~d����}��6M���Xŕm�ԳYa_)�G��Z��!��� bi�����3�9�j���nH;���/��c%fWo�t�B��P�z�	4ڴ���M��C|�t�l\��q�����P���k>��h.P��O��U%A�f_y�N �����.�B�b�E�׿��M������8������P�O�r��eY3� �"�ȳ�����+@תݍ�-�
b���b8��a'-�B�!���q%�����R�	�/�k��d׆3.K"�8O��4�~�=)�o��=�N�ԁe�XQ�Y�:�D������ښ�3 X>qOķ�OE��
�(r
�O&I�l�r�ȶ>Q�hz5�#�ļI} �C��:�� 3u��8u�]��УSJW/0}��ߓ�7��Hi�zt�St婿ǜ����t�l�	�rw����!(�yn��o4�8;P��[R���d������C�!��'MՌWd��D�|u$��s��C�L詒jd��H���e�;��Ѝ(�3|w �@�Z.tP���K�"8��p�}3�iJR��7/���q
0�a�l��%���I+%��V��l��sz��)I����6������Y$���!�1���s�/�l��f ����79y?�Xi�����_�Tr�T1�����#���(6�}hk���O�URZ��O�I�I�ib�E/��7jWK7M�C70GA���0��L�>���2�%��&�s�����5�"W��q��#��<�5�ұ*�?-�S��O.����
����l�-p��A~D�	�Z��''�u4��"�E�8P�B�sr-�f|BⰪS��
hH��ȢYU#J�R���w��"�N�Io���L,�M��of57�.=��h5mSe��#tڃ�edעA�����,{���M�XB|m{�y<9�v^Og��K�Tc��� �[ӛ�>B�C&�/%�S��i>}����|��s5~�H�F\B	���x�%�T
�VQ����[ 8�j�f$�ς��<�Ё�u�n��~���B���"e�J�Su�D���^�����=�ч�$��\�ϱ��+�U�l4���²�$�M��B�HaS�����ybD9*p;9��ny�N�J��n]զn(Нb\��9��ao	�V�3;!��}�����j�y��q�.:�kYqp?�~�����mJ�(A��T��^�����:��	.��'C����Gt�h�չs��K�͏�)Zt��okr��/s6Uv`����d)�>�S^�^��oCS��c�R�M����?���UF̎p�	V�!�+�{��?���Mڀ��_=*�I;!��Q��ǧ��}�s����HP+��k`�~˝X}m��]*?�>	�xцJ�h&����R��Z����i.1�=�n1�@���P�5'Q����f��9s&y֔�&�`����94���A`d�u�`�:�y�'�*�`O�+Mb}A9�Q#+ ��,�8wqn�2��B�5S8�n'e]�pq��#���K������bɀ�����y�����z����=�)�7\<;N���!�#Y��˾PA�&��fv�
�4��X
/�٠mVL�+``уy��O��&N(�\U4��c����TX"�}�Κ����'kqc� K^uoJίѶ1��]h*�O���t�	k�ްL�A��Ѐw����&���o�� ���*� B�WK
"*����:�l}������X��������i�<O
�s����� �fQwq�m�^Ƞ��NE�{�z�v��_�Ԛx���<��[���+�A�x'�Y��NKSv'�"�H��c���zJ$(�{'W��Ү�J��k��7��yȃ�6iT=[�{�[��İ��{S��T�0m�+NHz�^��f�s��װ�g��:*��e���= X;g�NW����fx�Ȭ8�
#�ק�PO�v�R?;݂��3x��^I������u���.�V��z2O���O_�K�	Q<7S^�B�K�1o����8�<L����VI�-�`4DG��������e뇃����i
59�_�듄A0u:�2�Q����8���rZ�X�VPGٍ��w3�-7�ۆJYj�������A�%�'��] ?��no�����>:  �}V�w�׸`��6����u��X�w~No�\��Qͯs��}� �?g�MB&�́�D,5fs�+ ,^>������һmj~���-��T�E��G����yX>.�B�W>�@g�yQ�ӵC�l\��\V�& ���c��d�%�~�M�F���Y=o�Ⱥ��(����������zA(	.it�
�(@>�ꥲs��$ 0ǥ7(.�I����:e-5��%���g�m{Yƻ~!�s*MB>L�Q�4��nf/��f�)�tL�V!���J/�ά����Wl"��(jȞ�� j�b2.�*:�-J��	��(��­��z�C��Yw�1?n������}�$��:�}�r�i/�U�6�\�G���n
�[i�9�������9�܊�T �tTe<��*��mk��
%�2���x��Ɍ�y��!t!zWz��]9�A���r�u�ؽ$,��q�j�	�9���A0'"������2��:6K�U��LK����'�'�dΐ̠�^5��wA�L�x�rY
Q���8���6�u���(�;K���D=�Nbs85��Q4'g���B��Pjd^���܆8�ܑp.u<\HRY㉸������ЮǔE��[�M�h��ݥU|��M�@�q�w!)�F�6��{^�O�>�³$�+���%��A�%��H�I�F�[���>V�x�}��)���m�C��l39�������Q�s�nH�S;� 1$�b��VFS8L�9�T�F�f�R4>}����!��Ȗ7��)M�� �{�W@aO���ؔS��`�=+�\�ՠ� �\8u}���W�8~�;�g��w+�y��5�V<y�=	�LD��"��c��{qF{6A���`RX-%P��@��������U�2vJ���^��0TAs�:Ͼ����h�<�z3�EU�"�ǳ��ߡFBQ�eNU� L���J�,z�P�CX��eL�&�W��N�/����f���t�]!j�F7�R\b��4ҷ��2�uV���JY�4��I��N�!�΀ˆ�C)��@�����7��>��F�3������xFW�DX/�"@;0v��c��/���tĽa��ک���H6�ڊ�J}����Лv�DP-f�����D�!��s}�-3�7�R�������������p]U�9���*��;KR	��kƎ�ja^P���n�f 6m]7^��e12�07tID�G�F'�2�w?zF�o�4�݌�:�A[NO<Z���|�_ZƼ�;dq�X�z-F�gJp[ܴ���ߵ�c�G�_$�]�X�{�<�'�� ��mv�A��ZM>j�Z�x��g�M���u-𯛿�Ң�*��V�����0����,JA�5?:�Q;ǦT#몖���H#$Y^�@��I��7-�f[u�5��/���@��(�m�^�v		�����Av�~n`P���n��bhz��;�ٲ�=�x�3�b]��Ʀ�"W�pe�����M�B���2�hr��Q�_��9/~Si�}2H�G���5�Z/���t;��1�p/�j�{�]������	՗Pot�q��YS�9��	%	���,�ĵj����۫��I"��R��C��� 9���v�i7y�2�3t��z]�_ҹ�I�"��+��Z�=�(�y����$ð���_싧�R�s��جT��g��^՗�o	iY�X�;��ÿ�h����2m,y��Anb��6O1�����n�=N���И��$�i�)s�g�S�7�X
�[G(���ڿ�`6�ǫ�r�eJ�@�+g�^s��*���{?���T-�Z��,�.��Ոb�U�.�
���x��������%G�q���M����qUo�d��d3�+Х�ݪ����T��/��|� ����;�����5V�3:1A�Ds+���J<h��RB��P	�P��DbAKVs�[���
��U�3|T�?��o[6�V�O,����a���Fֻ���/�t�#�������V�0�a���*tr�cK�� =�fڿ��aK�k�AV�3�r�����~ܽ���� �l2E�y: �L&��B)���a�.�QZ��$�䆸
�����~��J�fo�/`aQV�v1(R����qQ,N-H�Z�寲X�<��aΑ������69�b ��^ȏg�l����v��;�?z۾��G����oAa������5�[�ݹ�G���%��	3���8��Q��;�[��N[�V)�>{M�Hy��[��D�@��4r�y�p�t1HEn�>"nL��vO+C��5Q<(����6Nҥ�~������<\�Ln �+gVWJ�ԴT�P2[\��(;�i�>��<󗆯�a�g���xnW�T�E8W��]R�U\��L����z��C��෌�H2VN��8b��Ǥ�S�k{���R���/==��L�g���1���mN�����'��q؅y�-�	�H�/w{�P�3���
����U�� ����V``�*%����n,(�k�!1����>u"Q�s7�b㳹�� S��oX�3I� *pN�}V�zá@��ow�S$�����t�U�c,(�]�H��fmg4�nq P��s�?�|)�<C��jiN�sIێ����u�oQa��V���ǷWg
GjFP�+W���ݟ�NJ��ē���ٙ�b�<�)����0oX[��o���^o�
�N3�� Z�] gUW�����	��D>(&��.�2�n=fv�0�ۮ
'xΈ��dw�5c]�S�3cz��h�Nl_�hH�A���:�?F��U��r��Ǚ�#��\�ꗀ���l<,�w)�����
"���h@Aka�OY/K�Ya�K�ț-9�r>�N�E�*�F�X�4[��}�O��/O��fJ�B�=E��z)�򽓓��/����"_z��4e�Lg�Ӛ�G�ŗ-��eBz�Z�Z�j���
�B������Ԅ����u�.��I������W�I�p(̇��+�%)X%6�W�Vܧ䛢Hz�M{���냛8nȖ�I���עy��Wf��*<\U³aQ�~̈zHvP�)�����I\F���\*��O�p�6G��s���i9�m�����a���cC��A{�;��`ўn|I�������.��y��+�
? �g3�(vX+7ZJeu� �����{q���羫�'[��}#��'$	?�u�AW)x��ڦ�o���9���u�Q�Ll����*��./_s�;ȏ6���cÍ�8s	�9���j�4d�����2mL�
�S��s����~����u�n�6.UW�%�����F�����NmQɐ���Ka�ӣ�'[��������YY{V$�d\k�v����&6K��y�������d�J��1W��	kSn�R_�=\>�j��#8�`_ZKT���G�}'�����t�X��j<�FP�_�i1x ?3����J�.<눏��0j6�d��둥V{n��w��0�>)�J�w��+̩��C!���6�-o����@��]�K�o���f�M���8�ɬ�J�R@im�H5�c�F�c���MƩ�@�~x=̳�Q}����7���,����J�~���4����5�_�\�O{j���=,7/@�FXȫ`IA�$�$��]�U1&w���O�k���1w`�~Z��S����`��5Q�1�pg
e�����,��{ъqp�����-;r^���$8]^�{["�ڴ�B�B�ԈGo�gX}�ICf�P+Tu�'�̾�)�j4�`�l�w]~,�+N��,_hP��5῭=}�!������l�׃�8MQ��q�H��)��>-]��k��C�\f� �s��d��IK�F�Z��yi_ �X5R����*l���b ����Y��&];
aވR���f����娊M�!�1������:�#�eF�
������[O���A���F���{ 7W���h0(�Z`��S��p���ߋ;j��w4E��~8�ڈ��C)�����1�#4:h��ʳRR�p��n[���B�L%������,�Mg��Ӥ
�L\�[�l9(vJU�����u�5�1ǟ]��8��mpx�����~Nws�P*� ���b��!%�/�dx�͸�Ӂ/C:w\[��h�������(=����,�j�s���������gPی�$��Rk��>��o6��y��ɗ]Z���$� N&���u��MuԌgH#q�f}/<�����_�N��������A� Z�J��p�|mA�м�x�A�w@(w>��ݾđ�&�*$m�C��e/a߼��x�s�#=�⋰G�7 Y�>F}���"�؈�y�#����JVG�l�.f��kY�JL��#�/.R㾰~�]'��̙����E�x���?�w7|��q����\�e�����=�����/�����p.�t:�'͝(��[;l�d	K�1� �}��&��E�Ty.{�&�R������3h/C'=�B�y)СC�A1Ӓ`��:�{�nwh+K.[{����,�\|G [�v1]yb|�YҌ���hgGG3���J�|�rn�p����u�cݡ�)=���7�~+5\���5?���4��y��G���VS��	��S�Wە�9��إY�Q��6i(���R��
p��p6�.�A��l�*kH+�+�ƅ�pݹ�M%���l+ȧT9Q�"^���@έM!�AMi�3;��a]�|"�ڨ���%�,ڤQ������WĪ�cڍ��2�,��U�O��-*V��qq������SIV��z�5�6#5-V��C���>��u�����?f�;J̝�/fX�yt�����37T�w���t��*�%��y�$$/�!r�Lx�1*K-k�`T���A�n��G�A'��]���u�.���R�`j�Xs5��&����vA�`�7lm��AAztU���̉������f7
!%�f�
b7-�H�\������O�J_���$Jl�����a����\��N鸐���8��Y�9E��^�l�䦔�?L�[���
#h�[�g��*h?Bf�@R�6���������q�#�%�Lbt�I�)���"Kz��;���`��n��S+oi]�+.���^��U8��q<�¬�~W�c!����}%]`����x���39O���f_ �lM���ڿ�e�X:Ê�\�����"�����{6�%��RN9^��u�\U�����J��٬��Ǻ�Fp�&=0h'�Bq��q�)fN����y�m��Y˃��<&�a>����&ݎDD5C��Q���� �S��p⃏F�&��	�*�3\��V�C^�q�,�y� r��ӭ��X�4�}���8r|(���f�Ξ5D�(]�Yu��Å�^4סsRq���TPBm\ՠnõj��>��t�	5PO)�QA�Q����!�M�FF�/d��yjx=��6�z��9U���ߪ697(,g�!�Ɠ�.���tG�Ȯ�t<)�͇y�J!�L$:b
�D����8.���nm��>�i�a���x�|�x����������;Ǳ�q��Ǖ��1��"������bF/	/�>�[lM�а��P� � ��R���.0N�X�aw���Չv-�/ۄ������3�v�tմ6Ü ����K?F�#h,|pj�o���X��N����={�(��u��w9��?5z���X��>����i���i�AE
�Z��%\��ݥ����iv��K����ͿC�,�L�&Vd�I.�h�-�ǯ҈�1�r���B�~��C�b����^œ��^���{`@�kzչ��:+�|�RQB��:h�j�hcn|U�؁����tI��'I��Gd�6}��8f���eU��M�ىݼ0��������	P���w<��h-]�Q��vq �~i(%C�1M�LR�HT�s����u��� {<�Λ�q������.Lq�V�g�5 gz��������[tB[P�1xsC=2z���נ�m��qY����p���y6�:��`������89"f5�}�Lk��P����r�Q��_L�O8��<Ds�]%D0��j�>���"����� �"�Q�V�����/N���0;~����q/:�����q���@�dy�`�n)���F�L�]�铨F��e�Jj|~^~j��6�#���� ��}l�ܫ���G1�	�D1X���it�'AB��V�I�����hk'9!-o�d��(�m=�	 � ���U�VZ_��'��V�ƨ�W����a���f��M�<L�+��ΓPOJ����m��������sO׶�O����,<"�hb���9��B�H.�$qn��^U��Q����^c��������� �2��:�A&��b�ט��c��r��==�}WxCl.c����nKV%�����ƍ߮s�?�ڀ:V���Oޙ+ƨ�fj�1��sQ�O�r�{��T$�!q�g�17+�? 
ޭ��q�L`�H/0B�+N7����~��
������x�>!4s�qMQa��^�i�V
9Yr�}�����������>����D՟ּr<M�]��&�b]͟l�	,e�g�k�'���*��
v�_����p$wӌ.�������t�`�G�?�mI����x��ϧ��Ⱥn�B7pn�9FU��2t��1�@M�6�lh��_�;ާ�W�W����>��-����!2�`2�ޒ���~r ��c�b;'v����K]�3�Y��<�̮A�`�x~]�5�b�h$��@�Sv3(�?�$cP�U�_ �����y��p�Z�p�u��P���'Œ1�|E�0�3Aʭ����!�����>IPZ9c����=)"�MĈ1��"Uِdq�Zva�hgQ��`Z��}�2��b."�����fi����0�8َ��:��dYD_9E�vը��q�`����I�^���o�IiO�5�����0I�{��/�.�����~����_�Tr�V��Z�E�ӓL���WK���|L�TYO�\扐=��@�an�n��kW-���Nk8�)i����j��/�Wx�Gk��]pѬ��=����₮}� ����#`rG���u��'�2���]q��<B�f6�	ҍ���@7����fr�6�i��n�_Y���ֿ�SI�Lh^͖b�း�">�x<zx��Ϛ.�n��\��Ѧ0qY�S�}���gz%��B�+�w�f|ʝҘ�n��m8EL�0�]t&E~���黍����:㛤ÂRN��Д O\�buH8Q�� ��Wa(8��>a�����g��UI��i���� 8%���l���#ዩ9P��e�oܬ��U��g��aY�'wlS�N����w,�,|i��m���8�T����K�Lt����(��%41���,\��\r.{�A|#��;%z3�|M��G�$<�&&<E]o�����[��@MaZ��xB�bVB ��q���^����Bw�����t(��_�$�� ��}�M^��:2~h�I^	6��t��5r���k�ջ�P�|L�V>���Q�%cȪ*��~�6�Nj���k����	d�2{�k�8����Ɗ�1m�MU�K��qkN*���Y�����e������q�٩P�Vy�3#�HP�$'��S-�5v���M�T�9p����p����c��i�c-cq4�>��}s�ځZ�f��z�҅�Mˈ*͋���E�G����zv�Q���-����M�T��e��C�ik�*1�����L��3ҞY�
�{0}��x�k�M�Џ��M`)Y�BшE�)U�\��Г:�c�,f���&.�j����<*���1�J�������������%G��J}k�
`��L�;xkS�=m*�t_��>~!�1|��O��]��#�Й�:��ݢ��0������1��?�e��x��˴rv1��.�)<���u�<��Ys���[0���S�]��)�;.�a1�wp�\���+ V��ކ�E�2�y����>֕���V���YH�ϣuL��!�"A�[E����g��O�	�c�x�q�����\m�h�J��{8p��(Q�4GUL�C����-��"?�h��!���*O�U3��n�[��f]a(< �̤����ĸ���mKuSE�5�e�����R|` �̠��NL볜�>�d!��0����]X#���e���QLN�"<�����Q&:����/�� ��`�~m��9/��lrv�»ކ۰�?��-B�U�{��j�~�T~\;��q��(,�e����%�Ǡ�2��w7	s8z�|�3;*�b�@���`Ѝrz��(�p�+I��=W��ph3�?�M�R��5�E�{}<d�[[&M<%S��(b�	c"�i�������lct2l��0�4�uv��K�;��@ػ�ܣK2�����y��&�kEH�V$!�)�~���'!�\)5�ߑ(V9�,K֭�.�+�|�NA��y��q+�(eEo����tƛ#'�?_��6�בE2��_��+�Zr�S�q}������"X���%�-H[�;����o�7��Ta��Z�q���c�c߻�� �Y�	j�����=�G&�'�|��?�վ��J�T�
j3�A�y�=�H����O��7.���P����׋�������7ʯ���[����%�D^_5U�)�����p:{.1
s��2�P�+��]���	������Xo������� $�J�����$`2`�C�v>
�pN�X|l� �3��": +?h@�|�̟G"����I"kC���4~��1��B���q�]�l8m�C�G�Q<宋�E�����\���t��K��
�M)��{6���ݟ�@|
x�)a�Hm���4�<&6��4��g�;Ԁntt~~�f��#n@wb�;˗dg���~���.��&�O�᫲�!ģT�5�B����q���!g�r�KN�ֲG���3�Xjݑ��Nc��Юh��n��c�6��5���iK�z5�Dށt�l���"�����6�^�_�}cN�7 eİ�ލhY����v�m�%�?ԇTف��ɛ�����X��[���e�Sd5�����L�I��s���'c���T6/e�sefD�$�x���-X^���7��V�5Cչm@�z~�������@ʿ�^�\9+�_3��������W#�z
x=2�r(���k�.C"�	]�W�,a�J{�4��'��R&d���M���8+���eɍp(�!��~��-s6Y����f�����%���,.y1����Ijj����d��|������d �=`©?�Oz���"����ה��?�WݸӸ�P���<#���xZƑe��ӳ�1j<��+
K^	>�-:��*�n����	���4�X��n[�*�ֽ.jj��g-3K$8�	2<��0�k�ܞn���%�n�Bb(V���o�Ƽ@�>��AH�������[2w2��Ed&�}���&��r�{y�O�g��Ϙ����XI�n�e�KZ�p���pmY��[^�
6���t;1�U��mkt��d!�X����
1x'e�g�>��ws@ą�t�>Y�9O�;p��J=�RU_�,"v�`� ��)XD�~*Y��_r\��:��*1jC�����)�Z��d������k�-����Ӗ_v��F�<Je�z4�,��}��ly�%]c�A�ܾ*TY�-���\mW���#�H�{1P	J����_�����¦�U.���ነ�����V/�{[,�����Q����k�S�Ϟ-����I[[�К�Z�%~鄠�g��g˥�KMZv�T��jv��߈(�]j
ZL/���r�(r��
�2E�BWb�PRL�\��ؐ���?�]�1�_�Ԥ+�����G���F�� �QT�N��mv�b5zjb_�<��&ʆ$h����B�!�����tL6�YIY�\a�W���h�3���T�vUi���D�kg�(�tE444^w����\>g �F)y�֖Fўԯ��q?˛��
�(���r��_�֏(JRFH����(��ɧ� ���G	��G4���,�Pq�>l�47���b�
c'&�D> _5b�_�R\嫝ǌ�DӮ��io
j�BSˍc�us�2��o��wg2��=����h�Z���+����EH�-�DP�uA�Wa��́B�?�u�e���7!�~Y��&�������ϯ&Y�T����v�H$"͎��n��	У�;���P��a������SM�Sb&��ue&(E����RP&�-��f=0���Jǘ z4�'8~�8��]et�e�ʗ�l;ȉ��47��l'�1�J�:D�`�ƣU^�>"��d�x�Fg���ϊ��d u�9�q�}Œ�w~Fࡌ��ȒʘV��$Ey�
[6tn���E�-X:��w�O�aS"��>�M����@����}����&�a��v�P?����t]�<�@w� ��}Htu�G�V]#=?���� �=�{I�F�� ,=~�d�;Gf�b�B�Ŏ����C-��([yc��^>�����q{�*cfN��G��c׊�,�
�N�,�9Bxq�U�$b��5�6�T*L���>��B2]�-���U���@�Ty�D^!$y�U��Y���"�TFBi~�+��Q�6<�_j��>,����+�d��\_9��H�ś��TS��_�gw� �ɷ.����o�N�;Z���P��v�������.�ۀ7���Dc��"�	�g\
kQv06�-
	k���PJ/��Da #%�=�Rg-��J��������٥:��['�@��$���A0�J˳"v#�����%����- �_�1�ǚ�� Z:��RgK���!��2�X��#�!*����7������RG7�\���W'LJ΋W��=Kn��*f(������.O^�sW�5�wq�����s�!��%j� Y�t�'��d��<�E��o���c�<�n7/h���Ц7�湤ך�O���C�u�\-���~ۆE@��?��tkUQur�8�1v�Gz!I�������"_�{��B��p�S��'L�yI۰�T���/�!��<N=Tk�P�b���X�R0^�<�x0�� W���m�B���\��&��3�ޑ@x�nG��C�g��:��{0�-	z���Q}��3I�/K�>������U�֯�t�3yt���������(�cMc�T�鞛��S��,�G&#��sL<>�hO�v�6���<����=�b�ƘU�8c>Ba�1�:)��m)x"�	1����'�B�H9��0|S�����Fh�d���d h[v:68����C�R�W����n�}(l�qڳSN��xB�Lk
拦(R -\�G�W6%�'Vh�+d��a�X������7t�rx����"�gFU��_�(k����r�Zf�}�ք��	cO��t�囯O���<Ԇu���)�?��Zy�69����������,1��F�����:�@��.E�j�qp��}ڶ*J,�M�j�^%��+��!��	�������Z,�OV���e�C�݉�j���M�s��O����SP�r���N��ޗŠdD0QZ�ٞ��=n|�gf  �JУ2]��G�����:�T�z�-�J0�M8����&�®�����`<�`tٗ6�k'�������Q̽�X/����ܚ�Ç�H���
�G5��\�� ��pgq��8�K�1�С������U����͇=у�~��X�Ƿ�����Io�w��ٻNYy��?�ir��N�$�������\ek� ��1gXBՐ%6X'z�C7]P����������*mW>�$�{	{�+�(�7v��+��q/s����B�Mo7�_������,��GD�����.���A�c6.��gk\�����DI�@;Pf,V�˄����g�U:��?R\�p>&�����q��]�<*�03#��7���T\(��@Fqbi���Ӄ�X��B]`�T��V��m�|ʸ_�� φ:�hr.D�}ݲ�����s���;�l~=���tQ�J Mm(p�S�zu��7��I�ʍL��8S�p���i4ET}�:%a��m�J~]���~��,l��aa/T�jL��`�����_J��^��qje�0+s�a�q����%J�y��0��ia& �x��D�v&GVx����+e:#y�Ճ�酭��n�,�
j,.$a��3�	��-�JT�զ
��������k"��|̫Ϣ^��lc�:įt�(*�Yj��i�f:Oc12Qt��&4�����FY��}���Mb%pn��U�3�-��Æ�3���2����6�� �}�z���e��_�����CpX��Ai��}m�D�U�j�"=�Ce���O��T9qLU���.;ӗ�����$=B������fk&t<|A�.���4<��������	�=��C��CB%���w��[�`
|��h*lX����S�<e�_sqv,R��\���ZT�(V@����ϲos,�i,A��@SEs�)�6�ޱ����0�kV��Y-������t~��o�5�̾`���QKy^Pc��E�t	Q��n�w�* �ڌ�Ѳ�?�1d�?��:/��
A�e�t����m���@+��H!`!���˪t�4<�:�u���J��14l��.'�#7��	�=7 4# 7����pO�I��#��ѩ�E_�Є����ٺ7��3�i�iR��3�U
���������jmp	����
~X/s$��;����_
��6�M�j�!3S��r\((�g�Wt�����M����`9*5�j��E�0��t28`��A��n�d�����/����h�~���0Gy
��/bp6'�y���ೣ|�xm^}ML�s��\�C;�./���C�U���w�S(���t"�
�3 �',b����Ɏ�����KqC��p�V�+� d��p�@�O��
Z��"��Z�z0�.��[զQ�$�a���������W�Q?ĐW4��{�Fb����܆�*�"�D=	.1$���I��V��4���m��TAp��U	�cEBM�~,D���� ��d���I幡$���-V!y�x	��c_X�
��&2;N؃};'K�V�d�X��\�ԯ��2���I�6H�b��Y*���tG�cQ߾��s�q�TO��J�e\ ��܊��=s@혃� ���=�^��,��0Jpu~�| }�-t�P��:a�>_8A�a��z�P�l����e�i�R���&G$��!һ/��W;���9��g�ٜ�����k�X��R|��]����-n�G��"h��%H2r`e�s�o4d�Z!g�~/�����g�;���lY��$o�qzX)_利��jޗ��j�#3�z�}�X�jﲏ��7ħp�q]I���sQ<��앨�e�J{�]jj�جpvi��h��LZ�."	�����Њo�k�h����-Y��S�w��F\�����ǎ�K�I`(���v����܎�cFZ$����k���;,�" 8����Ʃ�QTv9��id�ؽU(.��c���K���UsM6���mc�aZ�ʍ�섿5$W0���k����f��Cf�#��EN���
��T-.��~�<�6_n���pW�P����c
��[ڷ�|���q�x�k��/2��|�L4�u�q����y[o{&�H�B+��[ir�S��;p����x��f%;p����j����CN{_@zAW�À=A�t�|,��E]���q�Z��zxL�nE|]X�u�\d'|���s�Vv�5��W"r�>�Pķp�z<e�c�%��_��� /�F&m�ko���| m��,	~�69��D�芁��F�g��q�#�5R�s�F�!}�\���L��d���ZP��ɖ�/��|��'�Z�&��o�k���x`ٲo��/�(��˘�UYb�x=�I�fƱ���Q��>��jR|��H�!Mp7ކo�~+� ��e���]CM�sN���������V�U�>޾�y��*�3���OV�a�K�n�����kGx�i6����N�#F�W����;;��۲|�Ҵ�ۅ�/,�sU\[0�!S�������:u��R-SE����H*���1��Q�b�\;���gYqc�&V�ѕ���D`�7��z�t�*���|�IZ�\�?���>A���)6������V����Z���p ��ǩI2�u�|��E�H4=������k�|y�Ji�!��$Gu�w`��-�1���I��V��H@� z)��ώ��&Ϝz?��[��[5C������s�9#'o���8g1�5//�˩&z��m�	�	�a�+�S����w��G=�~��k�������#�r��K�}�s��C���s/�"k�p
䧱/F���*��J�� �0E��	2$Z���ɭ|�b'S$嶠��,� X���©\�qUH���5hz�~P�-�����t�geR���7��$�}[�ֱ�$��!h�3d��@E_6�0��A	|�d�!���o��o�k����+�`�Tz�����?6?ӡJ�7۷#�`���`��1_w�C"�3�<Őݲ3{w��SP��E�b�1n�Cpw�Ad�Ԑ)�R��� $�ы��:�	���������D���P�JR��zw5�TL���;)�BY�D�p�sAhm�OpZmt�-<~o�!��=k�4���g�ᏻ��Ok /��<%��#��Փs5-&��C����a@��*N�!Q����S�x"�����ۤ�C�,:��Ǚ���ϰ�˧%�T��OyL��$�A0\�٪���� �g4��հ,�����{c��n:� 'X��e�&�?��I
��AV扪�i�s�ܳ���Gj����D ῄQ؂��9���u��^�=+u�W���E�d;U�A׆�*{@�L�$LV_U}2���;jW�y�����S��B�c�� ��ID��Zn�aJ�l�j>Ԑ����� ���D#��x�6XdP�+�`$�D�l�!��9z1�-�q��Yd�{/u�|�g)-VK��2|e(�ͭ<�T���� ܮv�1<�꫻��T��y������V���7o5Wx	~�'a�屙Ȏ`��s�T�(a���� A��W.6�6�r�?q#m%0$��]��a�
�ʄ��2��(�'x
���Mt��m���l��c+�g
àX3��~�rΝ�ۮ�E�Z(J��񺮖DC'�p�7:_̀yiit��~`	Q0�͏`�0p���)2)	�?RO�6�ٵ0�r�r��b�E1t �9���B�d!�����:{���
�6]@�ÝN����D ����BsծR�Q�x��Q��]b/�����v����r �F �Ƿ���k3V&��,��8������i)���!M~CF@�pG�	NJ5W�����V��m��<g�PG�2��>�|��&˂HD��s����d� ��]>�����r��K�ӌ�V��E�WM�
w�VIi���1�4��=�䇿����j�%�4?a�x��Wi��>�':Z�X����7����哝p���)�i�\G�oU�Z/"��X��fY�9�p��b7Ds��c@r�vB��OJ(�ε������}��O���xH�ܻƐ. }����t~5q'ac�����U�$�ڿ�I�ߗ��
�J�N���hw����ld���JH�#n
�(,��py�hU��;Wq�I���e��L�p�<9E�	��W;丿	1Қ҂Yj���&��@G��2!��M>*OM�R;Ui��L)��d�>���]	�ߗ/_`�U%�D
��\�䰅�Z���=�]Oz.P���n��8�a}�=n����� ��nb�۹,�ut��թ��΁;]����˴�L����JQ���3<G�_��m��e�g7� �WQh�m�-H�)Õ�\n��T�~/f��=�؍�!Y�˃�6>��k��Mn�t�����S.�W�qnh��w���#��r�Ox<%E~���v`���Xh3�e�"�2[����=�O��IŃ�"?�Q�s���H��=�#�S����P���x�f�4���-��z�]X��i�HA�4O�%iu��e��D��;=���n�p^�����@b~
���6#!yy֨]ˬ<������:'�ͬ1�L�����4"����)�ޑ���@���'��a�rp4-E�Z�2o
�.��;�?	�z�����6���1j�NJQcQ9Յ&�^�y���(�ђ�.E1�9\�������<+,�ON��8Л�3�*�I=��?���\�u�A&�*�ŁE��'�n�J��|��;��W[eV9u�9yn��9�<���fTUk���p9�n��5kaȾ��:�ϻ���j5F+3��	#�*�Z���?���U��$��qv>���MI������E�r�=��I�|8��ρ���^�Ky!�ϳ�T 7O�io7DL@Cn��7�cd��1��78ʾ͟	&@m/+!��A̟ .�P��{�H��Pc~��H���i�\~�%�x�.>=M-Ò��1�ɻ	�S��Z�6���U1�"yAt���Ex���"�-8kz���}
�&&I]����UP;�?Ȉ�0���b-�j�uf�`/I�5z����9����'A��b��T��\��Nc��cFȖ�E��
g��Ly�<��JR}>)�\�?�|���d�p�4$�ʘ�a�}�he�v�0�!o��:��mPp���wCn��K}k�ϙ��Wǈ�>�2o9�Xdߓ���p��^��]D��{��@]9�LGĢ��ep#� �6>��g�xc�|*@Bl���f��Q獨�a�NޔX�g��iX޹���9mյ�׼""D4�b�,��\j\~\�}ިĆ@�]���w�jD�Tˉ�c��h1�HslP凳-s:e[��~����IfXҿ���hp��Eۏ��6�ʊ�{�'�=H�<�Y�".�ڦ�W6���/3�K�[�
z���ťO��ʺZ�w_�q��DU���k�
'���RTh���fH=�hM���g��>��5���S��¾[��|X��*�fF��Z�zw�j�CM"�.�pĽ?��	�#m���-QW��Ŧo��ա���Q�_H�������EEC�q�
��R�YӶ��1 0J$H|�{�}�q���S��#�b�y�y��b��&2�E�д�~}
���XR���\d�5t���9-:0����V���n�+W\k����]o����K
��e���m5�!�:z*��.ٯ6�P|/��c[���k�X����p��%`��h'�1�[�D+3X0qY)�T&���o�oC5�;��6L|�qU��㾜�e�P����v��Wԕ���s̳�Z����ͧTHu=v��x'lJ&�uv	���.��d�)��T�Y��'�a�Y�(ym��xq;Η
w>)���H}A�R��$�x\5f)㨙�>�@XA�w�ɰ�;qn�̛��r�~���M��=E7G?Iry���#U��W�D��A��^ϖ4���ώ�K��̥Jʭ�TW�C/>��� �� �&�Wa���qy�Be�}@U�n�D�3#��~2�&�E	������@�fM�.�m��p�mgWx�ezD1�M��1�.�vq����"@`�l8���![�S1��4�l/>�����	GD�^Ȋ��4ȶ�l���=�D�!��D1���Xӵ���N���q�OH�f"�wҦ�c���u��'#+`��k0�'�P�Z�\ӛ�97�dnBnm]��#`U�L	3���H�r^��H"��6��5�"�<�F?L#����%;hZ[QJ���=`K4r���A5v��%����R��H������2�|��c"�����1�TS,O�$�Cc�{qOwT�K����ێ�*�:K>1/J�K]�B?�|����:,���N��׋mݻ�#��Ȣ� ��2�)Uւ��
�lw�F���8+e�`��ӂ������X\�u�K�hKt�!f� xq	=���~?RX�WB8&���oӯl ��܀'����#�6�9����(��H�	��ȭ+`*n��#�r˫kV���P�a3���G���$����Æ�)i��^�Ɠ��ڊWo��?¹�SÍ�S%��%3��:���z���G�\��{:���b#�v'�[+3.t��]�r�	���f�R�B6��s�<q�9*��*fhK��i�8�T�������ۣ~M�&�_��.�|	Bl*�ͯӀ*��"���c,�p̜�)�dWʤ��7�z�F>�C������9s�f��=.�=��.*2QBe�]�1��>&81`Z�e��M=n��Ɔ����/n�1�����7�0D'���͑\Р�S�<_��&��}�ð��x���>�����h �*h~"�ݭa�"����:KY�@T��,޽�;iا�KUs��Jā��d��}(s�\Y5������f3�� ��+ZRz�%M����%p�Ka�x�p��y��cw'$��괘��ՠ7�O>2M˙����3�T6L���a��N�[��//�����AY*���7�L+��oY�h��p��/}�9.�j��s�_`W��Vz��@$y^3j���������Ԡ�9�V���pM���[`c
6`�����LE������D����"X�����8�fBX�Z� �r�KP�clS����S�o��#Sj�x2�eܳ��/��y�;�g��3�~kd�x*�k�Icӕ^���_�ج8��ovI�?�6�|G�,IמL�\Fj�O���Ø��� a�3|Y,��(ƥ��A��0��s�{S�뻻��T+�r�<s��PzR(o=2\�!E9P�l#��y9bZ�7��R~�(r�^�#0O6	Q3'M�~��F��[n�Y���	����B�8G`�28��z�7�'��53]W$[�Mk�}��F�f�/�1yf�����A�Ky�F��.�F��ML��@;�v�15rT%�r�,��c�'�Òa�	�E�/H���z���q�>�T��|FB��m�S��YC1����%yx�J���0O�{��pc���nO1{?'r}%*4�J��C��H˒4�VX6M�!h�dj�����A-�II��N뛆��(�v�(��/�$��0�:�++���=�������ۏ
�[�$/���O��:2a���@O%3�O${��:G�����4��1oD��÷�;�͆Ǭg1]�C�!�9᠌�] l�d�M�[�^ρcwؽ��D �a��� �n�VX�o���S)A�0E��<y!$Ή:^�T����d�P�%�N@v�T�ߕ<�D�ĝ[~ѻb������Q3���1�xO�A:��T��n4�ciw!�M�M�s7n�a�r�xx?�i�kA�/�ʦ^�P(�V���mf�������e�2��ܥ����7S�=1u���;Y���ygǦZ} T;~1)u�~�^'W<v^Z��\Mv��&�ޘ�W��QvK�:�_<g92"L���1R3�t��<���'lR<M��:w���y�u����AL1��]��h��q(^O�6�k��� ?F���S�#�����U��bu̊ƪUI����h���������)*��>+^D�3���6^͈��w�x2�&�3s�������l��4B�!�o)m��D���1pޏ�S���R���ɥ��\(�N�(�a�a�r
K�ǖʽ0O�bLMq�\Q@sC��7g2��z�e� hw�I�| 	+܆L�mÈ����5��'����Q��&E��0bv�\��_�&��!��������Ժk#YD�Ic�h��=^ek����yx���p5���Ӻ�:t[,Iy�u�5x3脜,��FUS�K�}�ιG�WULwͧ�=B�DN&�f	&������a)Fh��/�\����d�+RF������c�;�p�kh����?�������DR�'����]2���,��5X�+_�� ��Mm�*ΑMz��O����XxzT��p�������)9OеD�zĩ���4��nJ	k[;��\3au�;E@�x����1��v*R�T��\O�ށ�Čc�`L�h+Y�D�H<N��[�
�B�j�g�!� 1���BP2�AM{8��`_��:{ُ,Ґ�cN��k�M�D�o��
��M�'��c_�c����t���6d��NC����[���ޤ�@�8%��{ZQ�*m���q��Хj������Xc "T�X�*a1�÷*\S���DE���V~
_gpeN�u��ULe�0��(*���u�Z�n�Qz�$�D�����F$����&sQx$܅�6I#5?�Vi[�[��f٧�D��໦*R��R\�L�E��׎���Y*��+��鐸w��%`�)��_O i�#�G^oه���B�ւv�F0�&�����^�^���R�t�c"��2.�j�����W����
�Z����MSPW�I�D*�0���_:�:�0�Φ(lsz�[F�% Zh�rw&�8!0?��@V`��)�ȹ-;y� �ۻ�~EW�+���v��Z<s���<�e�R����uI?�;���ɫ�:,�	Ѫ�꧛1��O�/
���h�q���)�&�a�:+�|�Z���ue=1�.���y�h���7���T����r|����w�$��
���&��R07s![�����������Z��3&�5�I砱�v��fJ}��p�ΓSi^G��A_��os'i��?%�L�-W���Q��ż��!��^�_`8�V����|��TK�oZ���� ��Gw��v�>
��u���6����wY��E�����f�LrZ:Sj' ��<�N-�;}�EV�-���0�L�M�����to�;�>���pUA�΃1���/�K�'�o���c�G�xA�-�(Q@��6��A�ՉN3��~�p�cg��4����ֽ���GD��{��ނ��f�~�$P�n�['�7d���-~����J�g���5���Bu�@��í<m���&����fܕ��J���q�:��GaӤM3��(p��
ʛ\��l�3����P.X��31���Aq����Y��vq��z�2�Q`́D�ȉG?��Z�2C㇎!ԲL*ն�IԵ@�[��J>�#׌�J���'�&�Ħ�G�$9忐�RER�&l\|�]8�0d)�lK��WXe/)�U� c�?ׄF�d�f��L��w�[�>ut*�p��R׽�4'�> -�8Uq�������2&�����k�F����~��h8�.a�f��}�޿f��uK���뇹�/��I���J�����ni�OP�K��̒�w�Z<D��dI�% .��8w�өӶ?e�Q�v��g����C���|m�`
�n��;) �L��\~#���GS$Z[D�ET٦�P2��70��{��R�}x"��� ����j	��@��&,�Z��(;��!�F�#&d��y���{e󪯊F%�srB�k�0"��αn�A���:r�9B
f���:���s���ܮ�w�i�z�ӹ]n D�k�C��/�KfJ�:�H�6��g�|�WI���)>�I
��G���酪��a�3�"{� &�ʖ�E��7�4�Q��0ڙʮ��H},z	�G[�r��Z�������	�v>8�sHU e�T�_��:_pհ�R���?
���|��_���zW��("銔�gY1N~
�q�h�<�C�G�°�"���e����]�w��-���V�6O�p�w�]x$�LĒ<ay�u�:C���"|��G̔/�|��#�*5��s#N(V7Ps���Ĉ���D7=אx�7o="K�ZU%�f�:eC���A�������9#���Cl[U��y{�*�)�:O��j��/�Eϭ/D�~���~�j�g��kl�ș�.'&�0-(��-:u��)�߅C�d)������S�����CX�-Y�%y�X��2Ѻ0n��5͌"����XXQ�6tZ,��l��S<���M�jHQ��.w�5�&���Ii`����#}�N��.K�����K�j�^���D�͂\�����������P�֗Q��1r>( �Q��`�@�@����M��b�;3�������a)J�2�j�����*�v~F�����r��a*�0Y?G�6m�tҔ�?`\q�ȣ��_.:�Rg� Pξ�?�f���2���{����0 ƦU3����w7�8�� P'2�qBC�fϐ�Z����t�4���B�u+��=����Ϣ���a�^E�Es��ٛ��ͅ���㜽�v�a��G`�ۍ�Xq�����i�Kۤ�HM8�h�7Jocl���p�F%�½͍sR/��D�ԇ���|��#M���Π�V�M.뾂x�3NZI7RQ�h�������-���Gg�ngH� �D#�Nh�)�14��H��۽��i'o}��*�(_�y�{��+F"O0�yp����NǇ/�ݳ��~��U�?���yR�Yl<_ۃA�S_&`m�\�d�W���Ȩ��㉋cQ�dy7�Xk�ݍ��j
xc9�=5ˌ�r���^���0��]�g��X���;��+mA�[�c���YE���#/���ST�M,m��O�;�������?\x�T��`�����Y�U/�z��F��1�<+���:���M6QЎ��r�+�r8C_h�������Eƫܴ�T>�}���5�+�mrwzE���?���ejj��&n�?R�5!�䮏d~C;���� ��Z{���д;�dV���������x��Nױ�7�˾'oS�1R��WvK�5���P��)�	Nt
�������11�c:j�ER��\��Lˉ�G�i_GD��O�K���x~?�³6�Z���������!yi��dꍻ�]!T�;Ƿ`,x���r;���]B�p���5�5u�Q�Sq�ǁ��XRO�y�!6��A��5�$�� j��Q��A�zE\ߢ �b�T6�����끵;����* 9�������:R��i4R��ЂS��d{&8�B��F�Ҷ ��\�f�,^^�$m�sҬA����J�>��{����ԩ��Fl�$-`�-9�v�S��@KSE: i�^Y�e^�R�u5*���d��Z.^����q2�z�6lv��W��5�����o7�5�k�.hQ�[�i���/Ͷ��Ihڮ �blc�7��8�,�M�l]�n1�<A�|�p�ġ�C*jsP��2rg�s��ģ�@M�6L��á�8[��ڄ^7�"�D�r�g:s�:$����H��8�>�|6f��HU�W���W���oǷ��/Q��}�`a�@%���$��j����=��IiNBs4RzV��Ffk�'R��^�)q=lV�ۨ���;�(���>Lķ��};?~o���V�r�h�J����Y�z�Մ��-�ޯ����"�@��E�c8���-z��IG+N���մҜS�p,�՜\�@�g+�19��"�%jB�C�L�1^�m]���l5�i*
��~v��U�:m�#h�6��
c�f%�rT<�_�dyl�	�4'�1��4	��GI�����m�.m��ȶ�$ab
������ �P��}��p��D��j�#:t�a��m��ޯ���TI���ǳ��8�v �B�m_���CN6�I�̓�
ە�b|v���hP��¿֪W��Z�-7y��{�N���i1qތ�r&�_Z����G�.����S{.n�%������ˊ3��?�����˒���;C��<���7�W"��	�`5!&c/��m��M*��N�bg�;gmF��oeUεWFb֣�{|�X�!���[���̨�ML����I�8�JFIb�Lۍ�VZ'�,U1����s�+pb0���7��	��R��_��:��ɛ��W:m��GyuӅ�c�B�JԖ_S��^���T�g�g� Q5�En[�,��ހ�/���*�É���T�eF��B\�D7J��� 3�����Ȅ�%�Q؎=�X�J�c}j�@��%�&v��pF�3%b��
~�̛�A9:���1}T�F	\������$[�7�T�2��R��m��,7'�P�������%h�E�P��7��ֺ(�q9��<r��jؾ�S�D�����V�GSP �Ps�v���S��qNG]�{���R�C9os�;i���K��~��(o�)����YS��(6�3l��x[kI��1 �����KV�B��jN��d���Vu���d�&g�4�B�;ɋR"Q�`J����Җ�[���3.�ȥ+E��9EDe��ؚ=�Sj�cL��M� ̡@9�k���ţ���~�>�����,�{��S�?!M#����[g�d�>~�LQ)@�Z�'��%B��[⪫�N�C�("�Bҫ�EN�1-˗Y܌?`���� �>�Ȁy���F`�lD��W׾��ÏVq&e�Y���J局�2�RW�H�u���C=I��*�Wk^��� ����vR~̼)��8l�����&IY6^��#C���p1r�m"%�����|~��*�������Y/Qvm����ܳ�.�<y��.C`��5?��G�/ڪ�N����oBԒh��c[�
���e���׌%Q�YUzl��z�q�)�,y"B��׹�Cd�?kA��B Zr.�. gr,��e�>[��=-{���Z�x�j�}nk��|]U��kN�1g�O�ڴ����H753����7�W��,�xS��gP�WE�,:kVIa��n��3�`��j�x�f�Oct��� �Pl>�6���1J� �os��|��ǃ���Z��4-j69\�7��XFz����uPE;�{>)��%9gf��N�Esg]���(�E�\��\�ڊ��]�^�!�^�K�,��1,P�7.ډ�Ћ��
&�Ha�lBH�zS����6�n�̾"�ˈ,;�:BCd�x��w���!td��b��6.L��T�/�Z:9%��*�=O��5�:~����y��F��:��ź3��E���@L���:�!N039���軗=w	���l0ZkfZ�{�r���oM����3h݁UA��(Ͳ��B�
���
{k4���.)6���y�Dv0�P�c��C�#y�Vn��>N��9{��a����^��We`���������慛�VYv�qw��M�'2�M��u�qo��J���;V^R��`�Ik�&�"�㐿��e��o�	��nD��Q=��{HN$���'�;���f$=y3I��R|N����G����FZoi�b�Bǃ���'N��H0�r#]Qͩg������wPKrI��x�����_���A�_Mw��A�N6�勬�q��wygh^?b�R3��
�"?\�����c>�/0~u,����P�T�5�	}<����ݦ��2��	�q��_mÕ����|����,Z�uݦ�;j����\�Ûŧ�>����gM�L�.��ɂ_����%�\f}4?eW�c���^ۦ�Sr����Vf	IM;�
ӿ�U��,x����,��js5��!�Klܤ�&I)&y�?�+��J�.��?31w��P�)�ė5I��j��A��[��<鞆0�ˉ�[�6�@>�-5�
�5��~��bk����mY�x=V�p Օ�8���"[U���.��I���Lm+i��_������Lv&d�2���R�
M�`;s����x�ᾍ�p�`��ߏd+�0BI?`,�5��ї�֖�p㾹׺�.���7m�C�*]0�Mĸ����6��Z*���R���UP��L����~��%�����j����J���!�2e� �Z �̥�����ʊ̟�j8��C����XRd�+Xc(������3�}���/�[��ٲ�.HW:��8&5)Q+����aU�ǽ��0ߪ����#W�]�rY������{���tEW���-{��YCUte�|fw-����>��|2�1ݱ��������0�w>*O�����|k���.��a+�����W/F��ȵ�m	�H��O��Q�'o&�|]>)�T�Ms��&�:Vi��#^Sq�m�_����À����[�D@�A�bm��BF��P��܁�6ǳ��9�a!&�NH���[�4S�!�0����0�/*����o�)4<����i�K�'����"R��t�.���S����n�1���k�r������h�i�.۔
ƪ5�;o�� h�H��&Q�C��� W+���uҚSR��_र-Og��>~��U�����?�Cω8�	<d%���,�cEa�Y�Io}@��X4�F{\����>�2,�J���{�{��yٗc�`ɭV[P���^S*ȧ��������k�p�t����6D2I�j�E!x�4T}�w��M"�pNꍗ�N#ycşy� Bbxw���[��4T:���Ҷ^ë���
��LK��;�;*d�e�=����Y
� M���x��W,e�3��h-x�*>��F�S˰t�u� ��כ�Gݕ-�
F�]wt�U�#�TȦC�������qGz��vC��qLL�ps�T��~�Wsu���4�AZ�]�E#���4|@���T��e������W�T��梙�Y���kX����+��ש���X��4c{��R��E�B03��)��A�W���bZ:�$��V;�8k��q]#,QCk4��H�����A$�H��]R1wE�Rl��r���-f�[_8 ~F@n�teU�����������?�q��- -�FBr�eb�!-�H��2����M1 q�d�J2�)N[�����f��*�@0B���~���C��U�'
�Hl�_z�:ѫ��~��2���s�4�&����җD�[�?][˒�,���x+S3����!K����a�\ �
Jc�y��#��p��:�Į��������u�'�Ɠ��%�e����C����xv�����fF<����x��mx��k�d6#у/�
�P�$i��7�'��?�ϡ���.�����x>u�6��0��4�V�Ħ!��`F�� @!�㽳x���2	�1��Dw��ػ���BYk��O���_
&U�s�&Ա�?�`�f���y-ٲ@{Cn(�H�m�H�'�+�\&~�g�gX" t�x]Wn�r|ƩnR)�^�@��#���S���"��T�ܖp�[&�qʏ����~{����y!P�c�%��a�H�:y�_�WI[lyUq{e��x���C��:��S�z����׭�j@�iQa�^�s�d�FS�^��3:���6Z��x��%L�Ya�(>��:\�z�����y4��Fj�s)���G�Z5��q7��Lw���5��HL٥h;��YS�9)�߶1>�T6�H����y��%wC��樂+=���e�ʃ=I����BU
���ܳ
Ρ���4p����̦7�`�p�Q� �?to�%��K��	=�D�d1�C=O1p�����k�(%E��^���b���)�W�7���$�� 0()�~a��g:��߿�	��dX{��8
�R�15"�B%cOt6^&�h��noQW=��u�S!Z��b$�{��ah���I"P�����X;�'�X�����Ԡa�+Z�[L���,-��B�D��u�4)�]Q�́��:o��UBș
�M��|�n��b���9f��������3"��*��X�����X=d
{��Գ�Q����qы n'���#m\�47Yi����I�V��v����i]�;D	�)ZX/��-e�R�r���7@'��6;�������ɲv�8	�I��h��1C��4 �i���X��<���O10s�K~�1��Q2ƭB���y����Al/�;�፭
����� �.u!�6�'���2Se��P�F�YR`��~��F�lt]z������βeh�B����Ņ �D�90h�a�z�S�%�M#�E論D�����Wm*�w'����\��瞯m�v\
aLk������i�	;�������n9+���:��En6�8�pk%����_ȝb�D�1�
M<�'��:D�~��!��F,]Ր����@x���XQ6S��r�dY ��MF���T,K�b|���~��?y��}�M<\�f�e醋�2�D�,�y�
5Eb�����_�+�0����R�C��[a��Pܞ��;��>|��~Q+4�V��k� 9_D�8m�]������G����epoR��CTU���(�F'�[9漷*=����W]��l��u�莭���[����'��yɰ:�P�KTVd�l�٧kd:O��8�7�'��6L�B�;`ήn]re<וz�BT�t>5���*P}E~����O�����P�pX�#i�8�N:t������4�y�'q�a�L0�K�4r�-����,�'b��Yҳ�DPϕ.��^�8SELP�6V)a�0f�|��=gAU&F9ِ�8 ������L"md�|p-��Q?$���k��v�O7�K��]q��Ϣ��(Tܤ86O���a`�_.V�*O����T\$G�T}���ډ�3/�r�$��jz:[��*�"ɮ���Ե���)`�8&��������<4����/�l:<^��+n����O]jY-a���j���+T��rޅ ����y(�-�4 8m����[�E�ވ�:�����H{w�zJ�`w{NZ���l��������ҼW##���n��VE�}	e@&���ۊP1 k_8 �n"�7,��Yp��)���T��2���%A���\������P�������J��ǋ��U��M�@Z�kD���Mh̰�t~�U�u�t4���]�j(H�
�?�4<L��[e�(�#ț �L�D�ٝ1��@���@2�����Q�e|W�-)T���1:b��b�:p��j'���X
��,)�+;\�!IO(,�����z맳Y=��وjm���Z�_��D�$��ɟ��:^����sXɮw��gLZ��3��,�����n�l�LE:��h��3�<�.0���K3#
�x]�+���#ۮ�k9�6.�I�5�M����A�o��T�Z�Gz�B4�X5~�A���a��� ���a�iC�+�{�Y3$��#����R�к��d@�5#ڊ�n%��eIZ������z2��JJ3�PS�[��]��D���>�ܴR7t�ZY.��V�`̧(��z���u�@Oe=v��<�J�nq�����쳫�?{�5D��l8�N̴ͫ_tF;Tϴ]Ab�Y�w� 0���m�|M���(2s�5j=�#���S��_�>� I܌jc �����L��8�ӛ!�Br\�������lC7�v�c�Ƚ��7Ro��M���BDY/�`f�U=����l]����ѓm�{�֢6函�Q�_jq
n!�`�?��ĸk��2���ǹ�1��^�6���q<J��Tf��#��|W���i\/�����f�d��E�;ME�6������Fզ?Ư�����q̏��$;�9���]�)'�٦��%d�G�2gH���0���%��R��S�3�!�wEf8��B�2Ws��8�,�.G����-d�G �f�0�NUE*jt`c��=;�ے�b���t��qS���ǳ#��sح�TJ�������-�>���yB]�x`MdO<m5]�R����qc���,$��a��q�*��~C�f:��sB�3��}y�����b�n4
;O������M�'�kWϤv�Cc������ox���K�!��e�	���g�A�˫�=��xOƘ����%���6�/��:λl�kڢK�\�D���	>����@i�{����ڣb�Xw��v���{[� A@.À Z�� ����n4:�DV�f: awi�V��R�t�}�B��;�9�H;�3fT��%�q�gB���*9=j!���.m.� ۣ���XVg�hX�n��r7�`/m��";���PW�6����'da�C�8�"m��I�-6\E��0���w�3�]�QT'ׯ:�L-���$ ��6��+Q�{��>P�*��Uh�wGm�;�h
5%'�]*����|g/�p��;�a��d���z�Čڔ�)��}�
��-e\@H�T̏y�h���?�Un�r4̐@�`P8�pF��5��}�挈e�K�A��un3i-��[7Zr�v��@�J#���A˷);��I�_�v�ie�I�͖ЙDY�G@��s0׊�o����ڶ�jwQ���{q�~(^��>|� �� �Q�F�eTt�:a+�Lt�r��vrEk 1/�Hq�j�ƿ@N�R� �����1��S6(���Օ�.q�D�RB�Q4���nP�Y ���	�I*�|�����mp��'�?'@N������@��i4O�5�����=c$���H���@f��z����<����M<���w�Z]�J��{)��G�_0g�t�@��+��;��w3�D��"߂O�)�bN[����|ZR�D��i�����X��9{�Z2����	8	�K�)�W|k���8sz�����`���B�#0���_R�V\8E��$�Ì&Th�8�(2�?۝Jh*�Z�D���e�(��X�ɇ��z{��ʏU�O�Z
h�l�fG��yO���K���*P����X,/�2�Bt 9R�(ѫ=)���ڎ͛�rRh�g�o�BL�@�<��[�'h��9r��� �e���	w�A��%��tc�
x�k� �4�c�˝�����6��v��p�x�ׁ�-u>�id|�"��Z��	�~7��!TS�!k��m�C��ydD=JY��'d�ElI�E5g�����A�����xr0�*ڔ�����!2����%��M{ϗ�,б��O�JmV�6���֘�"+���°�����U�����D�����=��?��vr.�/%K��w� IO�i M���]j��w'!/i��8������^P�����gcy�-����o�{��[��q�q6���!W�׳�sY2w����ںk�r>��[u��T����'��41�������?�ڪ(��|y��fh_dq�hˀ��r � �נ75]1��=s�[uoX��\:l9�i�%��wD�fΆ�$�z��є��t��{�z���!{'��oy�f�	�iI�1�vr���W.��dC��簠_���t���Ӈ�T3K!���~��p�ܦ����&�>�n��q�����S���P�������Q�8��Z s��)���P]ѝ�a�L*]S�;����"u	*�RΪwo��|Rq��X�a�WM� �J$ntD�#i/�C�<�\��r���2���j�!�����3.eا�
{�O��C)����K��4j5 ][���0�Lkh�b���h��*u)te�?r�����O֌�d����,�fǵU ['�i>�U��يg���ڗ���G�o>����B����l��a_c[l_ɕDLۦ	��p�`z����8���S�U?�����Ekj�>�9�E��:�E�3rt�d �
�͠�>���:
���W8�w�4�+�+�Wc`1��ջ�>7��Ao�* ����iq �7�<���޺����I,����I�@0��~�����V�O�!j��'���5�n�R l`~�ḓ���-��SDp��3涟-�'V5$��	H�����bJ���	Z�Jb���,��M�:o���xx}#8�q���Id����k��W�v~�(�}���}��������g �
1��a<�J��9�|�ۊp���aQFi03-�@��� V�(N�0Cn`|��3�4u����BǌĝDO�8M�+W�h瞴ų��+Tǻ���e ���.���:9tO��X��ʱ�i�����1
����H��J")g��sl���/ٱ�bП��֯��A*�~�n��<�q74��OJ�ݷ�3�*a��@ir���ܲ��	��{�dM��P��S�[�����Ґ���s���!�O����j�mxn��r]�[�eZi�p�G��u������x��Jt�Q��"Q-��m��T �v��Mj.X�+�rr�&/����d=��~P�O���QwW$�H{@r��X���~0�,|{`��Iz��ˇ�݈�STؔ�@�O�ܳLd���F���h�Ah�'Z��q��9�/���<��I��U�$h2���7�v��<�<)j�p-���CX����6k�8�lj�!�ao�@,�*0Q&��f�ig,�,p�|�����yA$�Q�iYhߟ�^��n�j���$��n�Q�����jB����A��B�Ʊ�z�~���,-ɫ�U�,?�
��_��'Ӻ�8��������{�v�\��U��*C���#H���c)n���k2�b�T���zB�c��z�"K��r�AY���WZ�&�a���E�o'�����]J�����D`��RԈ�h��j#�i�T�Z���2�
T��iP|���p�8�{��cuwm/��p`cO;�6������o��w8C��Ҩ �ofq5����uN�\`�����}�K��O��iX� Y�3�c@rPn��n�s�����纍-Б���A��C�ܿ���D?z��ՠ6�������]hj�ϓ�>��w�͛m-��%���5�f?h�Z���/�_��q$������_,=Lџ\��x{�]O]��QI���f�����c	Y|`���-��E���U�r��qB��t��ĝ��0^OH��GT5 .���T�9��8÷�F���v���ԑ�������U��FR�L�_�ҵ���~ۃ4���Y��!���pt�A��dJU0���䅵r>U���<��nh����@�K���áQ#�Γ�Rʎ{�4Џ�hꖴ�*��=A(��ʷ�f�� [7qMo�K��6K�!��wá8b����Fn�!wq���Jg� B������2A�y���.� �V��&�)N��
��C��K�b��@i�5�@�LT$qj�8V��TM���TgN�Ʒ�(�k��DW�ݓ��MT\��K2B9l$���F�Ps�f� U�t��1����x�����jQM����i�m.r�(x��!κH�*�W�4�V.#��'QQ��63X�K��P
NJl��&�$	� ��x��`ט!�|��\�Xٹ� Y�s�x�z��̯R/�MҘ%3��z܋���P�Wf����8�\%�mLU�0�ѥ~���T�C�6̇�o��5%���TWL⟱D  ���h� ��6�E.z���b���GU|���^�*�k~�82\}��;����9�\ I�nP]�ި"� k������(\Σ�?۰�0>{�b�z�8u�%�J�SU}r�Z�|M�ٯ0�mY����c�+?%���X,���ɵp�S�*m̿�(xF�A�$�J������쿆���Ӓ3$����7f�)�tHw�i��n�w����Qd�N�z!�;kV�'c��#��MN��,��	�([�#���'M:9N��U��U�5{.�JS�Vܪ
󸚅�|	�-�������a�Cx�񔵪�>e����B�o��~�BFF> ��y�xQh���ҝ�eހe* �(R��PoX��v�����$z!9=�{�!����1,�ߛl��UW�/{���5���n�\ѹ��S:.%t�؇�����D*Ƨ�=�)3��$�	CB��P��d١A���c<bq{�x�]�K������y&��S!�-�����M`���-�5P!s�=�9�E'4{J�-%f��W� � ������z�std�5]���p㱷K��&,�9,q�V�R2��i���ĉ����Ar!ag�� p�n`P� s��X�N�gK��0i���a	�S�7ĩ;�fJH��x��_\�����'k[¾�~�dg���py3�WI9�ѽ..�YK�u8�DG���i"�RU�����t��1��I�rs����5��ݯo"���!��*)%i�\rc+�F�MJHN.˯6R�}�kl�:�8��靖�7�l0C�B�����#��-��5+��F��餆J�P2�X���V���MpN-]�(�ٙcҤ�74Kb�!OPZS�w����Q�)�'X(Hh��.�T�h�nr~��t{�L�R�/��LAe�wë��+}V�Q�H.`;����d_��Y��V+��$n�&�v�@�ߕ��Y/��wl��xJ��)EI���y�J�n�L�+w'e���fQqلG�Z�0��T`��鳁sV����qn6���<��)�}P���]�yv@�S�S��
i
e��{�p*R�$��W��*�F�8Z�=F��#����M��T��WL�g��o���2ZN�u!��'Zr͛�Ӎy�7\����A��O�ͽ���<��V�f^=���kХ�XU��5	��w$G��9V��w�+�2�1tWn@&bJ@V�l?����Z^��u���j���}?w�e���}���xpw��e��A�@\�l��`��屄��4��� �e�4�.���hx��ǧ�ۇ�P&�kD}�?8����L���!ް�IF�+�׾gQ��E�� *�%R�P4���D�[Xx]���'Κ)[�7������o9��-Y#z��(�
9��։�Dtԧz^�b���ݖSxx>OI&��`���@��[��s.�s^��Fng0ޥМh(�spLA��V������l���|����vG,S�/�
;9"{Í�_8�G!��n����h�S=��3�^Mb�M���C�Q���l�3��������|�Op����N`�ת~v�^5�f5���"dC�HdI"ېb���I 6vX��y!L��l"��� 14�Q�#�#�56giA�Q{�=��H�w�	�������� �#h'
rR�2H�DE�-��x����X6{��҂�2@��5�K���Rz��x���J�SQ��H�E�~�<&_:3��?lmx�n@t�{�xQ���T^zм�1� _H>Ø��x�[����!.��S��Q�M�����!��K�bi��٘�h@߷C���fYv��DB�C�Κc�2yf���-�U�usZ�˨0�]����|i�o�C�RE��6�[�)�K�1C�
�ؚ��8�����M^i��Pc���[S�_<�A���:^�I|�tu�  �$��b�rLI��-ݷz�o�:N����� �#�"(��G�|�[�}L�Q��?�fi�5�'Xz��S:�,�����~P+�`���4�P�TФ�eɫV�ᇛ�*�i���m8x���VQ�E�3�S�$E��G
�΀�[��2+!�ik��/�����d�齤�n.C<�{�p]y�kۄ2c�͍���@��C��܍8�>���j� UƄ\��B D�N��)k���2lR��bd`�:�f�c���G�jh�X��I�6E9��y(�=���W��,��<���EЇ�S0{ev���>��pªe��ɍ����W%#2|&�'��cS��J�o1H�i�2��Fƞq�1deU!ĳQ��"b�a�m>�?Y���xm�R�NL����l�d���'�=���������O5�{L���l?�b;6c��$��^�{uEp�ã)�cHk��  X�;'���U�<99s�҇-�����Zn�&�����4�[��k(�t��+mv�N\�c�݄ۃ�d��Qx�;�T��`%G:��4_Þaf%
��cw!y�L� y8��	�JG�!�x�����f{3�QR��*l��ZNah��o蒔tS�����.� #OT�B([X��Ya��z$�ٯ=��h.�:wxU�k����e��<0%��[��'͗�p.|����id!��m������$6�EG�Y��d�7{-G�Qf�ɨh�snIz�ZF��ߡ�4���қ=1�M���f!k0����q����5u�9�nr�T
���NZ��<��<�$7��q�~�	���f�aL������~�U4��8W�aҽ}*	�\,G����^=���|�<p{(�lĮ�B�#��6)�u��*��%+z�?Q�}מ�8O'�؝4�nc�y	�]���3�iȍ�>�-k`L�xP�X�۳(����ߧ[oÞ���=$���YwYz����� 
���P�v��Y'��˯K)_���0���g��Č<�w<�sP��� ��7��64`�%G䣈cp�I�rHt���D׎�{n���3v�$8���,�?�׷�����91P:��@����I2����N���u��-�R��-@�t�!0���>GlC.�dh�աn���>���?�z������Jo������9��95�d�9Ș�9])��U���f�t�?��s�* r��{h)
�P�R��l��~�l�*f�9`� W��{)`G8�dbWg4X�M���-�xΠ�QKχ.��9>!U�br�����a\�W~0�:��,��5����׀� ����5s{��R�៚ E���̒��� A�K�_3�
 b\zN�o���Փ�"��]�s�a]|cϳ���l��MQ�]��ps��ܥ�p5*�wxu��|x����5������ǿ��Y�,^��"7�o����Q�b������a�sj�[燑�B�� d�$ ��!��J�[���dNЮ�ҫ2��ߍ}�P �����vV�~.[��Ph�aZ����ژ���H(T�b���=`Ë(&)�˼B4C'�˳��AxC~�u�r]g�d�� -S6m���hLy�re; ���߹4������6"�a�dE�rgdP��a�m(��5�U8��,�8�:M�� m<͚�~�<��I��M�3�5k�h"���d��Oe��آd[w��* r֣/o)�tZ��>��X`oY��`7	�Z����;�a��[}�\�3s������"mJ_Ƌ�-�4�?�ali�r3\]�F��]��(��KyE�
�����bm���,��{����D�x٣+��NM�Ǔ���Z9�"&;" �߂� 	!@�:���G⤘��M5Y�l�=�9�ǈ?zc��Ɂ&��h�c*�DT	��F��/���������.o#��]^,Pi	G"��K�3��['w��6���@
M�U�	,x�2�*y_'�%��_���;3��9��,�uD���{k͉�/�w0S29��H��aٝ�(��x� �% J�0�s�F6k��k�M=7T �$��~��t�I�w���*@������=�Zh?��d�:���I&�2ܘ�{�(�cW��hf�I!�y���ju�����|?=�t
4��mH4Bscwـ �ZCT�J�S%d���S!9�dy��IE���ZU>X����v���� �"d����Х���}h�@���iwު��H0[ik\>h��n9C���r��X��-���:tj�$���$�S�ý�@����U*h��~����������e��8'�9���(�>YI��H���srCx�M�I�|lo�(wo��oQ뚶�+$ŨN��w"_�ʘ{&BU���q4��$r�JR������@(����ޔ���!��t+�>�����������+���3��H��%���l.�ntW{˼��tD�����Fw�T�6 |�]�\I�>Uǩ���f�Gns~y]^�+lT�����O?��I��o��k[h���)4-8�S@�C� ��	�R�3�-rM�
[0�/�&[&|�X�>g�U�>�Q�o�nT�LĶ��%MW�����r'����1`H?�~G��}������htQ����d�����EIuڋ�Q�	�����

n����C�n"T�k�e�l���,?6J*�]��8`���i���_�|_qq���zqgX�.�*�w��P=R�Fp�0�h�ݼ{�ҥ�1�ʚ��{4j�B�E�@n�/v��� ����8������@��ѵe]Xm���`>��*�a�G-����s�UD�/�S�XVX^����gA:�_��̿��&�N$�H"[��uj��B��ck�,�`]�i���@=����9�J|`$�Y��y,#�s&��P��AdȨ���[q>Z!N$hv1���j��Y����F���p�QG|4GCTGVu,�T`hD�u�'-�P�g06�ḛ�K��s�U<�Hy�z�-��֧\�5��}�ձHg�n�XO��|�k�<��o9��x��-x���3� �y/[,�2��VQ���а��B��p�}�ٲCƓ~Q;N6��*�`W�8*�V�V7R�"U6�-s31��� ��7�48+
Hϕ�$2Uq�P���Co�\\��Đ?/чWH1��K��R�lc��r�s���d봆�]	�d-up��zY��m4�0���'�`��;���+����qr�L� �l�Y��']@y�\�|](�ZxX4� �{��(�(U3K��(��@os.�O=�.�Xg7(��z֭�9C�� ��J�d��Q�R�▯um��
�H�Y�9́$G�W�]�KWs�o���
�䱙�A�^�P�ˊ^�S݅`J�x��8��!�^f�ݭ��/�*�Ň>�K��32%��{ĉ��ջ6���PUe`ԗ�`�	��"Z�a@�[���b-0w��/���<�b�?O�C�J�JO�q��.���͞{쫥!�����
��G�u�$�f#�>B�>_���Y��t@m��o��}�f"��[�py�k�_b��+č��V�AҏW��ʡ(����,�2m�9��K��c������{b}Z�yf���5+�'LX��D�hC�BnO>�������� H<��Я����D���]l��|�3�Q����@NTE��4*x(�97���<#����Bȡ;K���4����&{D��d���{���ް�k��?� ;>Ϳᇀ�"1�����gw�Aw<��`ir��V�%ÅE������R5����֤ �ĺ_6lUZԶ'�w+�E�Y�,-;�6a�y��$�섐(͙٭�Ĕr����F>�@A�LE8N`:<���T�ۡo7���6���7�׈ �썐�CR��fo;��L����BaO��]����6KB ML:����M�v^ݣ����$c�����8H��!�3�&��@���V�Q�,iY���H������h�Y�F����<�%iF��N��
q�� �p�wp��PI�z{`&nw@&�Q� 1g�a��(R��Mi��<�W*)�M�z��L{���vb�$]��Xa�A�r�6��ceI��,�z�gӗ�u��d˳.Q�ч��,� y�9,ܪ�����M��/O�����P�7;��َ�՝.�V���PY�S�D�h���߸����������Б�Β�CԑW���!��!��k���u�^�H�Q��=��\a�9e��.�d��7��=��ujr���¤Dz�2{K�q�4[z;}��02�`ۖQ&�a���_�X����/����_ �4 ���}=�Ol,�0>H���Ss�8g�6/O��)P��m�VZ�.��'�A�L�(e^���,�n	�`9rb�	���2��e6ėI�9/�*�QM��v�5�XXL��1�\�*�@����.6�蚝���Vj�7F�*cWcSBS��U�M�����4�q��a]�=Rdۺ��e�i����2��/����E]Ww�� *d�p��DV�Mn�Z{�'�N }a½��mW���Z=�����[+�{$���>�i��P�qN��gn�e�6C�y���ӫ�@|��t��E�hQ��A��]�5`a���!�s�Z$��R��=�6�!ׂ"Z���T2��E;��9�!p8��\�氥<;����-� �	ށ&D��4��ǿ�������-*���b�>�= �;>^Q�<�H�9pb��R#E�i�n\��CR�����)fs�����>��"���Y��a޶�7�����Vu�["�B����7N7q{�/�΀��Y�?:]�1h�xd3"����������҅Q�ɰ&�R�7���7�\Q67[n��g�*�[����v���Wm����-�-		��+~.�E��\�:��03����v�T`���Q�u�a�7��#�0,���z}���y��r=4P=R�LP��v�
�M�7�T1��@W��σʌy��}���Y��<��p7�kZ!�+xu��5J�7 �j��vi�B�Q�SciC��i��������"�8�r����i�o �Q*���������z���qJ5 �yB�w4���I��#�X�KΊ3FW4֑o���7�z�:�����h���g���x��J��L�����<�t��5g�3J���y�(k�^-F-��,��١4��Z��n`=��ͲOWzu[�U���C�&N|�y<e�����P��u�0VwD�u�<�%��ł���}&�6h' ��Y,�%�F&v}�2�����������j�����Xkz~bJ�0k(�yU昱<w����eͯ/�E�E3mXyJ
�/?d�	Ϥ��O�T�C����u�$������X%�;�yy���#�A�w,��TH���^sI��j�=;��Nⰰ罋[Ơ�5� =��3��[^����q���,���O`E���L����4��WG��5:�q��������L��l�R� 	���]�&�-@=�:T�X��<�("+��Si������*���ޮV,]���k��0�.zq}dvyQ!k�h,�/�����}l�ߟlH2+�DJ�f���	){i%ڭT!�g�|Γ8͜����SY�����+��A�*^͉��Sa l{��N��G������Sv�O���o���c��c��d�C�-2d�f�q���{�~��0T�tN���V�¦�[�����[}DQ;zD9���&��O$Ch�<�$o�gP|y��@�䁢>5���x�8�k�FSE]�փ�4�(��UN�-4(�.�ϝ�w�G���A��K��%��m&��Ɗ`;L��T�!���bS���qJ��1H�K���<a��:O���9RA-��;��]aRK��
W5�j(cE��O+�a�(�g:�t"w�k���^
����.&5o ����M��V6�Y�"���(
#�p��g�V' �&f�Kb)��Tʄ�Fѳ?_H���6V����ʏB����l��[���r�ζ�A��[=b�H�()��1x�toOv�\��|q�GJ��P? �3Z_�l�"=&��☂9��d}v��"��EZ�C��E�t��i�L(�}k��jS[y��օ@��%p%���?&����c]��SiM�B��ҭb�*��Їs�Y�<n�	��Q M��e�'K>eʷ����D�k9� �f�iA�F�!d	�*�&P��c�M�,��$��I@0��L?�_�4��o��FFF�.x�<�T��1��_�[������n�B�^Z{VߕctE=��vh�7^&]d�f=bH��(�'��-�J�e`�Pc���@��k�D�ZN5�f�ƒ��W�����]�!��u��JV#㨠f�>��n���S�Ky`�m��o�#�E!᬴�Dib�ds�4�v���>1�����h=)��w���Q]�/i�u�bZs}
,��Oݬڪ԰|��I�<�'�F��Xj�7P�JA�"�yo�aMR��R2��Sk���Jy����^+= xzl�C24�K]�_
j���������E�ˍy�Q"�N�I-��J&��� )�wܤ0�RԱ���'��U�K��Y������/暱H+ddr�\��97��>��Sg]��[7��v|o�S���c:p�"�k��
��5 R~��np/�����G^�䝇	d)w�0vo�r��]7� �T����o��M7g�d3�1Ϻ�[�q�>k峺9��@���[�u3�d��S7��ʁ�3f�?��a\����z�!�!l�?�ՅJ��c�����ڹ���5��T�+��^��R��#����/�i���t�z��h�Tf4�DpT� #� ���&i���f#	_y[o��¦�A3@���Q��l߳��5c+�>��n^�^Q*�u��
�cV��ߵj*���tb�"�{�E&��es���;s�;s�,I�x����;?�4-Q�.��f�?ܴ�M�M��^���w`�}���"�U�C����� &x�!�jVG�t���s�~�����9~9��`�0�F�B�����>�D2`h�}�&��>@� ��7H��`��)}k߲��HW寳=����Dp�
�-�l`�g�Sgߌא[��#������w�G��i���9֢��]��c�\��X�X̪�~���O�z̀'G��ӵ^XX�>��۹��τ�&B�"� �t�XH��	4���7�2�����	ȱ������p=����6=����
�����N�C�Nc}�`�}f�=�գ���#h���f�^mO�eHl�m�B&U�%S-յ(�ڌ���8�mb�gFI����vS�#	�3�w�C�"G�D�-���;X�՜7�N$���ȮKJ�E��g��f.�y�x��V:&�蚰�����_X lt���X�HP��s�߅6���58�����6��]t�
�a����f�泇g�g�p��;��D���	P7;(M���t�C��!����*�4�}������ʂ����_'�4���G���x9�)�O=ؔ*?F3� ^f&o7N��O��e[΂�%�� �s�B�x
Fp�X\�k�3��Ւ�#/R�V��ߴ��_��������A|�n�АЂ�?�EP�F�4����@��� _m�F)3�R�n��n�/���+�Q%��n���58���5M���b�}U"��n���Cgbiu\~�v���x]���I.���RR����&g����ӛ�Rs�;lù��5q(#�_�V�/\��ڇ�Px�N��.+��'�b{�D�U语�d|�E-w9���N�E�x]d�>S<v�k}��f:�%4�W�����P��D{��5|���@�����I��:����(�6��j�E�N��$��Ay|��5�f>�3򢱺>̟$�^���j��N�nj �sU_`UC���n_�����~p�X�a;֕�Da�U��9f���@[��P2�,�uE̗�_�ѷ���Q��to�EI���ؽ������U^�*0V�Yh&6�$�>3�]7P_�#V�c��1,��:��bp#�5V�u>�2(���b�'�p��/Kb�X�?���p9_>l��.�J�^��ҦV�Gl�M��~�����K���U-Y:��:mn����jn:7I��Oճ��ă�2��H$��}ҜY%	a�+��G�R*���,k@��u
*:�r���wй�xXQH����/�l��rK��b�P��� �>=i�<R�6�v۫B�j�I�	!cO��fµ��v	���yd��?�5�S1�T6jaI�<K*hs�8}���=�}h��dp\=F��
Ջ`�:��z���{SB����b \Y�z�y;����������J}�f��(�9�!��~����D�<j�R+p>XYj�ݵ�Ԥ�&/֌?�֭�d�#�cKO&871&K�Ó|�� ��E�k7$�B����{U����?!|�_�R-��M�}L0r���0\\b�k��fB�fA���am��)� �_�Pڕ�ڶ�A�粻�\��?Z�i1nb����<��,��W����f$~�3�%T��ȸ:o%y�My�AY��۟�����U|��zQ��m�QI�l��5��mh�5����91��$M��T$sf�ȋ��Ȼ��9�T��w`��^c!��{#�oq�����f�v��.���an�J�IUHv�Om���ȹ!aL��#Qo|,X+a��&fYҿ��n��b�)�Π	�T�� �{�rT�E��b�f�9?S*F�+lU�q+�R§Tb,���A�����x�Z� �w��c��u-/F����p����|
��m��@J�"�������q�5	��»�%a�O���>���	�������ʝ|�!�Q(���
��hU��Q��y��\�'�����0'��
���ܛ�g�(�h��! vΨ%�0��M7"��XK���=�^��kY>D��p�����"�Qʣ��ʘ���2!�,o�`��5���@���8_BG�JF�b���G�y���t���|-6��8(@r�{�Ԣ+ba�-�Ϯ�z��2X=�[o9`�7+}(�yE�S��%MP�Ay����v�
�Y}j[|ё�a�q�K�r8		���u�M!$G �IrE�#��� ���EtZG����`P��!�ô��?���;|Ԝ���\��;K9>����Ö��7{Qc����):p]�d���$���G7sŀu;�*�b1�zx��EeN
/�޶\���f�=�O.���q1�����џ~{�sA�E�r��sn\,����-�I肱#@1b��i(K�қx��<�R����ik���	��"������Y�;!�*vG�3��J�.E	
����ӑ�W��*J+W��E�pd"k��.?�8��N���z�dfe��~��k�� i/�����w���rk.ЊhtR�Ŭ������3�+�,�;"GP��9*�/}HL�c�+��q�7��rB�[���3��l�.����k�TY(� ԑ9����Z7��J��� [�-�8�#oJ�4<t�mk���@��w�7��v���D�\n�c#{G�K09���?�����ln}<v��N,�Yc~!ᗜa�by�Eԍ�	Ȋ��D�V+P��lW*8����1c��Sj�=�N5[�'�&�k��E\�jvUhz��O"��2?8��%�aZ|#�E��U�Ir��W�<��]����"i�S�8Y���-��۽O�/o�F�޻q1�-맘5~b@(��1�1��-�8�Z|@��e�~P�j���F��=�В�i�r���^��Il�c<��>��I�{غ�/k��M.���1�G����ao����6�v{_�@4"�6���a��-���՝W��?z��������76_\�9� �l8[s�o�T{������;0�E�o�q���\�Ğ�	�i$7z�#��E��a8����&��ʛ��;�XД��V����G,��k��SU�t�SK�{WR�R��x�4�zM@�A�E��EO���T1�uh��|:���{T���4����UeQ�t�߯Be
_��d>��XG[����m�T���,`�)��΋me�k�].ٗ�l�� �$ã�^r�w�����j��љ���t�04�}Z_��>]O��a|��{��[�dq�ѭ����oD4L�{��o�;D�!���	�هǅ
�H���1}F.u�bl��T�K7X��A̩m,��~��-ź��&�"9�{)Ǫ&��#�r���B�*��';����(΂�@R8������8n�[`�ӡ(	"W�GfB�*���$�L�V����X��^)�Yg��^uK(4��^�v���ď�O,�'!�ђKR�kf�����ɻ�էŐtbτ�'H�џ@�Q"�9Z1w�WvC�d�����lC�"atX���#@)�bYd�l^��(p�Α����6~�Ɇ��}r~���ǩ������|U��e�+��[6�=A�N�q�4I���Z����?��� @�5��&Ye*�ged�|z%��6��ݰ��Ȩzn_�󏞎�ӹWs=��Qz���qE7V��ӭ��ǹ?���r��A�n�%d3k��kʩN��\�MV��R�2�<��0(��#�-6���.��
`�W���Ha\(�gQh���5�H�y��WWIｍ�!�G̤���oԓ ����iR� � u���LΑ�;J����00=A�k���A-��X���N�'���Ꞣ뚃�i�x�l|����/�@���	4p~y\�H�G�EnE�
��ն|�Ί��lF��"bl��UX}��� �*Z�^Fw����DkY����1X�/�J��k;�Κ3»��}eE��$��y���4"#�8~8j%Z �Pe�*%i $��L�p���n��!������(�L� [�Io̫�z���*s;��/����&��7=�Ws��� �-��Bq�7q1�*KOX���ۭ��.��8L���͟�S��3&f�� �`8[����	��'<�=Q����q
X�ϥ���?��$��uS�OO�5��C1��A#"JKr����D� ᩎNV����E�7�Ldl%�a���\e�%W��'�I�9s���yڹ'������@,��ПKo�7�=niF�CS�(JA��$��l��}�g;��R �����&��vɯ�n�jÛ}Z$���N��hE�0��!��j$__��kF�ۭ�Kn� �`@"��vf��Ua�Q+5�!Xp_i,��|��v�5�Gl�-���)�x�H�U3�={/�(�,J�&�#S)�9�ݣ�r} z�Ё����DR��Y��S������6�#e֘�CrTץ���4��r��!	s��������	�+��\D�`�Vt�&��?��R_��<�)T����X�=	�9�<6��T�D~���cN1�L�1)i[�:��7@�!��CJ�U�1Lj���O$krQ���r�����1S��X���<��2^%S��3a-p�?�0�F���\�3��⁧��?Vx:�v'�{z!�o�1�����aN�6�'b�d������	��4�e/z
��s��e����{�P�&�H���!$�W	�@
�@�u��&��!x��`  �6@I�]�H�'�5d��2��N5�R��M��a�weH��e� �VFW)�=���I�A�@@O�B)�h[� ĝ���n���\&?wh���2}���A��0k(�i���JH��xM���$�{	g�G�!0����V��d��R��GƣC˰�_V�����N�=&�F�
%�����B���-�ӫ�/s���I�����":�9�T���}���oC�� 0���6Q|����V���z&	l5�6����i�'���I����u�&J�qv8��%k���Sn���<^��H5����W[���7��jXW�A\�yE�O�{Vw~v=%;�X��O�8�,MJ�����)(x���p�J���ݫ��e�/	���#� �C�H�ǂ�U�w���<P�!�?�E���q�1�v� suݎ���c����46�kR*\[��؂�� ?�]��x�_%�_[ͦ�iRL�� �^�3'�f�Y����*�Sу����l��:�x�X�Y���H�j'Zq��P22��=�O�!���]ի�[G@�}����L�C��=�`�!R�}�\��Y��kݰϿ�c�hW.�_�����`��=A���} �Z�� ���j�^x�X'c������4*�tF�7^��ii�"B�|���E�hJ��o��?�\�v�2ȅY�g�A���=]���DH�s��6�����]]��]�Y��d�P��pHչ�z��G�R������?%���^��͖�U���*�55��[JN�D���֛ TV�(�WSΈ��7B~�q5D_C�����A��f�M,x'���w]�s{�&���%��<@$�[�LF�g�z��IQ*����9l��r�,�<n��b�/�>����ݡf���9O�Z|@Q�=�b��:�J0���5@J5�@�h����%ĸJ$��M�{�G>N����*�`��&�P�q�-�f&��.1\�)M�B0t���O'I������Z��u�a�8*��*9���2Hq¹u����DgNa�V�2��ʤ�R7�l��0
�,�ڟ>1��ꤹ{�o��Y yq>-��w��\�b/�|��Nzϊ�J�����\u5P��Ǉ�������Ԏ4�S��8�gG�g��r�wq��LJ�zr/���%�H*O��J&6lR/%����[[.W ��n��.�Ր�)!����e����P��JKΉ�L�H�Z]���?8V4��l����Ħs�;Wg��F^�|�Y]y������ȧ�*D��%^�ZalR�ˇ��.:xOx�`I�	�������(���Vk{QFU�.W{���k�;-M,�}��~�|�
�-d��C ������������b� �u�[��Ⱦ�I�?�.��1p~ͨ&U&;��l5��h�m3�\Ҡ�&&ϫg,�Z�-��-9�4̮%<��5�T��H�h����V�=��o@
.ڑјߌ����+a��C��	�z:��/x �hF'MЦP��*�=��.�W�ޜ%B!�wǀ�Ś�]�V�b�RN������u*X�`$U]��=��$���e��]��q�Qɰu��Yn��%�%lW�Y���)�݈�������qn���K��AZ�{���aEl�LfD3Q���[�2hG�����J�|�f4Oe�u����yɀ�.^����I.Z������2��+:�qu�<8���+VN#�4��c� �;��A��-ې2d;�:�Ff{.���e�*�y �u�p���;�y{'�4���?:ep��Ș�L�v�.n*Sڪ:t�̐vX�e�1��p�*_bG
*��?��H��25����\
QZ�d�XtQ5�s/2�$3���f�G������R�En�Y'�9bzO��n��ꞡl"E�����X�V~7�_&H����I��n��Ϡ��o*�,�N�vVױ�g�ڽ�10�Y�0ͱ��1w쑣7�Пv��]b4�	�o�uy�y��
o.���u�؁TP���{��T�1���2x��/b�jʵ��{�-��g$H����^�*\ō-VH�9cpv1�R��MVW�KS�=� [W�0b�^FD���i`����P����eN�W�6�A��p�r"�ȉ��}�qGD_HKkK*�]ZY�*�[�|(QY��ɘ�s��*G�d�J�PW�RlQ
~�#)E)b��[��(���X�I��bo^��`�����TyIO�����bR���@��
iƪF�,g0(��09.��b�5RF<JƢ��<�3^r����h݅�%�L�'����k�3���GG�v�qE�Z�U[- ��0ӿN�"��"s9�es���M;���Ua���#���P����A׎I¨�0�Do��$�gAލQ�.�4�b`�>W��2c�����y./.��i�$�ls�R2;1^mޞұ���*��X�k!b9>`
)�9E4P�ھ�A姴TPELjO85
�C��%b�e�B��v1������l���[�<k����n���d����Ӗ��9f�������S Ԧ��C�c��W"Z�����ry�֫�7Z�d�˽	�`���p�� 
��1r�׿�9s����ɝ��;��,$a��XeT:ǖ6� ��G0�0ն}�p���*��v����~�M���{����h�cgӑ{��Ma��KdD���lR6�Pv�s�V�t��F�;��<�O$ل;z~o�2����!�e�� g�	Ԝ@�	�����:A(��z�ʖz���M��(l��\.���J/2xs�@�DV����C�5�1��Z+��4b�v�T�k��վ�%��:�ݻ_$�6�Q������6�4u�Õڂ,�_�� ��Z\���Y�t��1$�MTr�
���牋Qݎ6�?��<����Z��I�:�^���T �u�iG�n����z��,��~!t�1��+`�}c7���}�OHê�&�俌����t+L[l{γ�v��n�i
��U���T��҅���,sOf-�2h�����z�]��^��F2�����?Z��F:�¹�0����6X�d8��xxj���z�����Ni^���3hz�Y9�=e��K=E[:��z��;<��]rJ���}���~I�q\�}�L�|����`�<�k�x�o�}7W�D���o&$s��G�X�r��
��!z���~D�Ń�`yU^?T|�!b9﹡����K.=�:���#�u�Ӆ��I�K�n*�:��AY�(����U�o�Sb�W���q�G\B<�i���3�M��Q���h�N>G�����5T��D�l����7��"�}u׸�U�	*��v�\a�7�M��L�X%-�8��u�^����V!�@%x54n���V���-.^w��N��o��u�ńU�+�}@	�;Z��KU��g��J5}�Dȗsp��E���ϸwy,�����X)S�V�-J�8-�b&U�[��S[�pi�6���
���NA�=���w-P!X���S���^��,&�O���fP�@ԘW?�	(��	�r��')��@�&�Ȁ�-�x{Ip	����,G���� �����X�\@��w�߯Xz�	�<B^��_�n��$����Ҽ�e�}�l,�0�J�+b�o�eA���r�+Yf����FQ�;�K�;kM�=X�aT||D?��D�qpZ7����w��}{�e�ѓj��{T�s��F���F`���i�4d�':ċ�g��ba�W�K�봿�[��\[�u}�|���ӘsN���:�bSp�#�B�wv�Z���� `U<��f�\0�J�;��}�m�%/�H��=m\�9 �0��E���k�#��x�������2y�N�\��lGg&�@�Y3�Z��l�}��i�@��a��K����c
-�C2����c���V��K�N��fK�u��� ���8c5��X�߮�Iw���p��v�� ��&��;r��T,��&���yZ�� ��wc	E	
��h�@
Z0�!� ��弯%����KKjS�$�6�H���Ϫ�[����pgd��r�0��׭x7?~���ɔz]5E���Dj����Z��L�ZS '��c�Z�zo�P©+u�?߼�^ZB�<��a���7W~��(��9���I(��M�d
Cw�䥿��$B4h�����JZ���-x������V`0�A���,�u��	�U����F���P����q�f)ts��Uˬ]�˅W�e*���_5>Jݒ��%���P�Xc�S]�^�n�V!�M�,3v��z����$������]mm���h���!u6�:�̓>�gK�2�k��rvy��ʈ�� ]�eo����Ag��!��=����*��H{���8�t$���ܤ�GL��jFo�i=��L���D��ӷ5v�`���U�O���ĺ�L���D��Z��˺T�p#rx�_�O�A��3t�|��Tr���3{ۨ�Nj�7J�:������������[����p�,JR�ĽCK?D��!�~B�:U��!��6��.��,
�X������Nj��T6[�3KI	EΒ��f���<�\�%'����{�������~�	��Y:���E�&�+ʁ�����2�)\�?C"���������*��؏�-j�"BP=E�lG���@�ϒ�I�����w
Qb{��(�q9A%TN�o��ݳB����m�?�Fsdo�$4�*?(/������� ��ф>ugT�ʮJ��3�(�u����_�O�l�|G�Z�;�N���K�<��u�{K��k��p\�t���{o���b��;�eyy"����[�{OД��*���ˉ�������MӨ��p�e0��ݗK�wD��ⵍ5�j���O�X��y�ݭfd:�T���9�f�N^3��g�����������DoC�v��n�����}r�lK�Ԩ
��D����f��97���K�_�����p�4RJ��\�Aм���]`�`-(�r���kԐ��!�Cw��'�@Zt�Qs��9q���Z|R��`{���K��i9���Z�H��ep:-�2b
��f��0	�7��T�ϴH��bz#R�W��I��< ��`��a&kpA�*,����	��b�O�&��[=�K��_.�~�P���D�|x��<G�B5Gh��ј!� �����@c�%���/�7��6��D��}�>� ��71�;����hE=>9̘l�k�Y����J�V�!-��	�̣R�˙W�v?�&������eė�d�G-)��@Mz��O� �3��X���/�[Ϥ�<ƾe�uWv��NX�v�׺����i\��Zl��f]��|}����(��=�c�bpU�I7a�^\Fw�TU}z9e�L]4,���I"�i�ù^�V��Aj�����Z�יY����4�K>iU��?G��9T�US(���&O����� �R�c�2w�͏aA�c%��A#u퇭=C��@���rd�}���2"��ު�S7�S�X��� �Y������)S�n+�Є.���^  *E�9��޶��ˬ'��k�ﵨ!���) �+��]O(�Q7T�
��禮��y�5�=�u��X�8�;�N�M�#T�V	S�N9�6�E��	���b�,a^>Ґ��Y�S����02�!��P���)K+��Yq��f�g[|/{�B=�ҮJf����50���s�{/���E�+�s��M���q��O�6��C�<q�_��Q�;��E�i��P���I�W�K�@�t�	�����n���?#<#v��Y�������c׮%�< ZrF��#4�XO�B[��^��E��П�Y�S�'��@�δ����&��VkY��]\�٢���W0��c"��� K�j�
%P��VΣ��|�J^�o���^���"5e7�"�\^�{��y�Ε�o�~,{ы��C)�[KP��
9dg�uT4U�2Ε
@����qE�a,�ף�����1���
f��
��i�f}���i�B���C��ӯ�7)�@ȳ������$���é���t���ӔV脹��Ei����/
Y�k���ik�xC~!�+��\��>�N~�f� t*R�2�K�^
:6'`�|�����agH�6.t�5i�W����((��:&�,�E��i*�.�*�\�؛>i���z�>ꔿg;D�{#�z�Ky��� ��]C8H_�S���K5�?���Y�B�y�V*]��!*�5�N��6�D�����Ek@�.ߪ-��^�܊ ��Y���/x�P��
b�H�ZdO<��6��βq���z}Tq{�t=ʗt�4i>��r���|��AXM���	�}�85��^��2�c�2c�����Ebgl>
�Lׯs�Gr���bi�] eG��Z�s�� ��hG�I��шeU��a�ϑ��!5�F�9���� ���9k%ΙL�ꀝ�ID>�
��b�?���]�Jn-{� �(�8�1=E�z�ēr	-������ю��|c02�+*D����A_�`|����!A��D׊)x!�k-��F#?Z#��Փ;���"F9�j��ܜdv�<I�ӗ,M	#!O���ES�V��іU�1�)>q���%ފv��*-���L��o��r��LV�Z��ay�r�݇��Ǐu��<�M�B�fZs�!�A�o��bx������X�|
3���Iu��hG֯�����`��?��x��|��P��T�}n������ߏ�0�����敯1ڋ���6��N�����
����G�Q�zG�gRE��X�'R7r������+�VT�3���24�9)���.45�yd��1���]z�H-N1j�,�S9�~�\H��x;��$t���ye>�[�p�f�z� dw��	'dӧ�6�bQC��m',	Qd�C�^�_ �Et�k�jJ�8�魣��W(���,8��,I�b�-���h<ۙ~��^bE��ȹ1�d�u��/X�� ���5���ւ��C�����6�0�����a<)���ރXFC�>�4�晙�prk$�D��
�.-z���|=���������@jw�bv��Ql ���!y��iD~p�q��廗G&�ߋǁ겓Xk��� ��2������%�T^Ԇn��
��NQ�A����(��^߮�*��*�V���o�z�q�!�V�Շ㟈�4��b#�cI�&��Y�Sl���gB��<��"�|��|ԐKU��K*�}�
�݁Ȳ�ִ�"&a����SyZJS�sdP�H�_���ї9o}���n���t�F��i��~$��0�K�̫����q��Tx�Szj��0��PplcCT��rl_1]�=C�<�}��i�"�9�;��!y�N��{?�(��FW֔^D�挾��!�a�ُ�W��� k���g�K�L��:�6a�Ǝ&���
g��^�����!����:�=y�/!g<����k�k���hgbz&nl�"ϕF<uFd����&�҇��޾��g�h�y���>b
g��k�t��'X�r*ܿ�9��?�\��Iw��Z�	ݍ�Hx�{�ƕ��ê�.ǭ���ʪ��D��.����E�\�f��9n�V�{v�F��~0��/l��i�$��P25��Ӕ����������!��5�yֶ�����l���xB�}��L#�P��wN�9HTƌ-���Q�-_tW1�3�H��6�����ګ1b�G��&N0�N�>��T7� �6��	���1k���?���M�%�A]?��٫�X����lW�M����?��gu:��K]�q��3�u��`���z`�Ĺ$f�(��.��MϪ�Dl o���I��}Y7�j�8���)��`8�E�-��H.��3IW��� �`��&���k���fF�X�š�΋��R�]��e���xI5�E��1Iۥ���<��~g�S%�P0/�U�����ͳR#V��^����x먹̢�: �$����P(ɸ�-�Yx����҆��R�|<w6��0Ise{vᶶ������o����G����W|�f�2X &�#��Id�TY���f�)�O~�>���,��m�a�-y����S��*	{�d;g��eN�u��&��0Jo��0`�Gi�����YH�H9�>�U}��L�Ja�5N�T?�쁦!��|L�R�?�(�
G(<j��ZIEt?�Qi���cd
4�{�(�E0	!9��&>�w%kM�Đc#H�	�¬�j-�$6���ú�:.b�LMJ��x��CE.�x��L��Ӛ=5�eƓ�vov�������0t'�$������x1$�l�W���e"�����L.�oHcs M�OS�b��%�]��`�����b��=��p��n1����"ո{���׎�P��ȥ}ebO��PCv���΅ʦ� .�0í��_M�Cmo� �u�
^�����ѓF�Aŝq�DA������^��d�~�͎�f)#*U�mu8P7[5�vj�b�>�n���H|y�Fڷ-i�Ԭ�:��:s�,�`���=3���8��.�Ul����"��a ��3h�˥\�ա�����7Y����F��Z�@|j�D���6bk�ó�� 8�ؘ(@@��H&�':�k�a�V�xl� �^֛�>�D �����g0��]�h���J�lz��(��˂C�zCdc���jl��ٱ��4�ﶿ\BZ�u4�[���p����0s����-e(�J�s{x��=����"�Qi��� "�a@嚸�#�wA�S���(���Ì�Jǔۑ�6plR1S��[,�N�ǯ'p��A�����>�e�+T:rj("����	ȋ�혋�5�-�J�M2`o��iEV���������yS�%����dbsL��S�?�O��[�6Ty�\�y	�ym�,����kί5Y{D\q�X������­����G*__֞�.�)��ßO�}��D�ʋaUze�u"��eEHV�ُ��נ]�v.�^��+:�~����U����{�)�ɛ��Mڐ눟�̱Z+�������z�IB������8��|�F#���\]��)�Tf���z �3}�\|v��h�f��0��6�[��ױ�����~:�pt��W'�҄r�@�E7$؎~v��4�f~�U�-���WX���]���a5*����HQ$W�d����h.K����E%��v��]�����C1�]�f���r,2����"�i�o��k�^K�z��Y�{��`(r�t���}�u��Ej^�]�;SB0�mh�d^DPL�觃:���n���,�'�z�
�.C�����S�f�ǵ��u�QY�����M�:3

5��_��r��_��ު w)�d:\a����/;y��I?��
�� ����F�ة�	�w>�8OA����6��X�%�ù��zA��O�B%S��ϗ!n�
��X�8[���T~I}<� �(v1*Q́۷q,>�T,k�e����=��Cm
�dڑ�C}+r����Ejp�zB.G�=q�]I��M���������?�5�6�М��MN�E1�:�l ��w���L�П����̩��A��w{�ge��@����6�n�Ġ���k�79�s�}T��0uw������2N)7f���#�sj�DSZ��)�V�f��a�]�q�)������PA������L�-��3�o�0�����r��Pp-�g=}4�v�����\;�u%_����\9`��Zއ1�o��tq>:,)�c�p5�GEf�?��1b�60�C*L����DbԌ��.�gԲ!�d[�]0㻯L�7����_]�6��n�n�.�	���ϖ��	��`�"q����h����L��غ�e\�n2�;W?�/�X�|�V���i�=C}���{��oJ�Yl���q���82+5�amE� ���Ifl	͢@�--��-L���������2���t�ZFK&ʐL�TۣȦ�ݐ�`��'j~�z}�=l�0�h-{I?P� 6����o$M^(J�2��k+�12�)�횇�
ҫ!��-�����z#�;��;BQI�f"t�X��%���j�\��WGQ�=��E	3t�����BPi��ƈ�[Ϛ�+��؝[�ێ���G���
�췇��?�V��z`�j�&�T�:O)���K��?v��c���F5�h�CU�~268s�E�2l�� yi\�Y�KA��U�!b���Uhk�('j�ө7�/ì�B�p)+�x1N3�ȔE���|{�b���RVN��;�gK{�<��k��� 3f�dNS�M結W'�������(9�1jN��'lj�%hS-��7����*��<mk��[��w�ͮE��I5��i}+�C�=DI��l���,�K�g6���V��}/�凩�A.�=�}����2/o=���_W !:��5�3X��S=5=X$f8���]� C����A��:��ݧ��F�"B�O/V������wZ�n@�n�T�j�o~������h���Ĵ<���gh�Ѕ|E���=��?��S v�Qo5$wP=��0�/��v��0�D8"g��z~�[�ƒZV)˧�I�rx�pO�;��g����2(�u4aQ2���f�)���5oM���6�/���Ai�B!�	9�.����R	��m��}JK��I�}���z���ޕ�jo�="]Ր\C���#�D5��t�}�P�@��ݟa��F�YP>�}��2emZ���A�K�,��k�V�g$G˓Z�j�{e4��Xi�m������!������;UY�kat��#D�믘�|&��٤(h���Im�����8����2���K������̝-����������-cd��$4�u{�:Q�`{	>~��֤�������%x>�KqO`߻��{� ��> 
x�{���d,��+E��"��aޟ^�U����ۅ7�T~�XQTƺ=�1;�Ɨ[D&;��Ct�
�̔��Nl�^#��٧����$j�'�����0�RM�r"J�4|�#j֡���E��{��3x:�"��5��D�X�ia�*R�j�ֽ��:J#{�����T��%�}WūN�����L�.��ʈh8��߹�C[���&C�j _�m�A0�5���D~�0yW�����%����$� ����ʸ�!�Ў����J�T�%N�>��f����T,.��8�5���6p9��-a�
�ܥ,��D)�v���gX��T/��"g��6�[����3)���?�ڌZW�+�1Mû�V��Y�����H�Hd���{ȳV �E��[���?l����i*��$��;����T��r}k����~!����H��'��T����i S��(J�w�5��=�;+��Ga�YZf���j����A�%�/���(��oaVuu�p�o�**+���n��9���7���5�.^��R~�
��=��#
d�H[6 )Y�p�[�v\˄�����g��x���bv�b����P��b��-�{r�/�����.��cfn��Q���bs�GYK<ׁ�T�+� Yu�|`Y���w����2��.r�u�y��w"`���˰v>a'���F�p6Ã���# R�c-��JA�c�e�$)�u��V�:K��O�)�S��~�[ �ReG1�( f%��<#r̿���@-Ŋ�ع�FjŢ��-$�:ߒ���Z{6�A	9�}Q(��6X�C6>W-���*a)\KѧȲ9���H���!Z �����#�hs,�{>:�T&N��z�.��N����q�/�mB�"�ӊ�d��02�E*��Y,��!V׃�A'N]b4���.f��+ߟ�����d�i�oS����� �].Фz��A�kW� �jH����Q�V�0��y�`��6&��@w��)͡ЄS�p�V�Be�L�M��u�vԆ���Ŗ]���H)1��������f�ڢmAw>��h<�
�۝�4k�k�墅����2KA�� �_DȊiͭ1OQW��͵<P~��@���0̞���]/�Hh�'
�C��Z�A܉x����7 �V���e��>cأ�)�:��i���b�� Өٝ��E�{:jh��� ,m�DrPS��!a~|�Ev��m�#��Wa��Ur��M݁�ƨDL��CFm!�J[h��Z�g�޼3�-�9�8�k�`������3m���D,�w�R�p�)Yɻ��\ǟ96*�aJ%�c�v��}7�0'�ݍI-{��`�춀mO���^�S� rڑ���}U�a�Q�+"���}%f�d�'ڑ��uD�*�flXboa'�!��΍^�lb���]Jsv�MT�6��+&\�c�)I��@Fu'=��]ʗ �R�5-���H�'K7o�ػ�^�l�<���P	��߸����_e�n����J~�!�1JE6�k���Θc�Jqa�R@Q�^}�1�	�B$�ZD:y�FI��@l���wۅRY���m��bu��0�8!������b�5�\k�8�a�\�>W��8A�N"^|45���}םa?��}�d��D�tjk�޲����N�����1�-y;d��ͮ?-��sA�(h��S/�)�iq�/A �(�p���$��}���hE �\1�9e�A��!J��L­6��(��ڙ��T}�/9���x/x��Z�x?����[
�i����%�����#�ܢ� =<!Ei���4�������;Tː��8F�{�4''��̋$F��<2D[��٩��#s�֌+S�p�I��s�c�vU�o�U��B/^6�ƼT;�n�V��rK���:fW�����k�wӥA�l#M�X��Ƒ�|����4�V�j�l��h$��!ŀЀ[�1��J�L9�?�m.Agi4���p�L��-��9��1����}��4J��� &�S���$^p|/s�;��u1�;޾$U%;eC�JQ�N�[	��M�זZٖ�߆�?�R�1&���� �;���!�D�(i �/���։��X�WUEu?z�,���%����,"It�xt��^R~��[�p"A�$����j�N2�&?����s�%�l"��̓(ސe=��ݗU��Z!�]�^+�y+��+���4���a��d!&UY�ړj�wݥO��sV��]����̱h�����g7��a]	����I��$��������K�7nVC��'sn\��_p���P$�רw�,e��׺ctb-�D�������FWw�_�|#���*������D���[2:��L�z���Z�eO��[�JiF>\�� QT%:���{�G�D�蓞%�� _���i&�@�Q�C;k�|��J�f�g^����3�p�+@������NZ<h��]�IV7�t7�P R��l��>�� &�"��/���T��[�t���"�vQ�� �rZ�9�ςŦG^IL�C���$V������HH����¦,��N��,���qy��̧Ρ��?T��T��:h�CH����V%nQ�R�P����2���e��#d�9S�>6�S�mn-W`�?nJW7��15J������
�wi�z�r6�/j�`�R�qp�췓4#3�D9T��҅�u��	�"led;3n(��j�%��� �z�->���|7G��r;��0ll:�q��v{~����CxI��Ȅ���g�X�����nO+Bѵ��1O���IO^9�V;͆ϝ����(�#��	m���Q��E�N[��U���/�L��E�Ƕ�JߖlE�6G�t$��#gD�@�s��j�1�#���h}�	����7���p/�g^��{�מ���A���E��F �'QmѶ�Zn��	ao�t�X��pl���h��V�'���]�Z�K���y=�s�����Y���w��w�LSU!�'rDRd��ƀ���J��h3uI��װ,1�?�xol.	�S��8C~Ͻ�<�k�9��s=}�I	(�#�_�ٛO�H���}֡ {�}	:g'v�|���;g:�͑r%�q/N�z�W/68I(Ő�N6^���!�b�R8غOҥ>
����aS�0A������OWPF����7��3 �׈�N�Л�:�qՊ�����љ?�>)k����?���?B� I�����&��T���B�g<�:G�~r��#r�6���$|F�O0ʽ�����Jք@��7��9�Z9�Q���cru�j��"��G��ӝ�}p%$�>r��8�-���Q6��?O4���$F�	p:�Q%"��w���V��{�w9������u$;qeS� �_F�xkY=k�ʮ�j�yv�Nw��a��ⵓs��թ81�����Gv����d�Ɛ�A/pz�,���lm��(�S��x��[+�	6 *��3Vh�Œϛ��Ug}| ���L��C�9�$��Y����ъ�r˲��Q�_�6?K섄�
�<�_���g�xQ	)�ᮒU�����%ݞ��6nA"?��F�Sy �����e}��2�hOܣ�i��#;a�+��N�9ǌjF*��H��hx��&_��U��Ĥ��q��ޜ�{ȗ!�a䗿D�^�߅�RYi����?��,J)��x�iN�Pj7�_���8[ө�,3��3�Z�T���W6�� z6�*%��
t@dʜ�4����(R�4� 9q<-}bHJ�u�u�:��J����'��]h/y�j�����U�]������8j=hJ���i��%���s�\d*��K�RZ�"'G0����وS���g+��;]��NR�[zx+��L���~�+c���P���a[ ��ܨ��g H�|�����,�\m$�p Nhc�)v/�$��4|˓����4.=���)c_���Q܂�(���ٛ�"������'�d���[�.� ڃ�%����E��XH��TE�+3`Ap�~���	�I��̕t�1U��8�����T<D�[@��6I^0�S�^���Q"���;�1�-��w%�5�e��v[����[+(N�C�N� �x�.�|)NCg��H��7J\U7��U�����H�e�(я�Tf��|�%Ou|����`Yn"�ʔ��&U֡ME_�2hDȃ���8E�̕�w:M(�RdA��vTl�V�V�<��� �\MYW,7�9Szy�Fx��١w$�Ӎs��L{�$>;{4!G����#�f :3z;�v���Iδ6�L�d�k>GR#x��]�+����v��_ ��b"g�����}��bo�8AH���:�X\�L��.u���a�ܶl�m��m?	C��r;��F����^;����q�I���[������.\
��9`~Iw�����[��`CG���a��,��4bh7����c"eR�-
w�;�cJ�Q�����i��
h$̎�!��)��S��G5B����\I���JC1�˚�9��͢Uo���~�c��X�����q�C�|A�g#ů�Iz�%g��!�V�H���4�P�K3��_���kj�`��C/>Kw��vqS����#��ːF�Z^���5�O�eJl��1�h{���ג(,\A�fcaQw`��U�?�Nǆ5PEah��Eږ�x��u�����?������የ�U86����cƷt��B(��cz���ޝS��a�6F�$�� w���o2�%���@��j�H���g⾷�f����vI(P�=�4� ��y��p�]g_r��Hh�@N9���G5y�,��	ek"={��%�x�>.��Bv�o���Z��g�f�����|�鉦<i����GGZ d8PFB���i{����;���o��k�2i�����k�������������V���G ���7��{{�B�c�kg�u]�J��bz�^���5I�~��d/��O��H�aI�]B#2w��]p_���f08�.@����	3�8<�rڙ)hT�.J�2�k��k��Pz�J�7
H�	D�A�������X�W���ĕ^һ�B�0��\���(�\��m��Iq�8>�t�G+� ń��3TRZ�t7�"m�,�Ҏؒѩe%I�o�<<X>��6��mu��H�6��T��w?@�Ơ���1tT����j�%$��v��H=�3?IB��/9K��ΒM^Q^�î���$��Vgt�|����G�3��P��}�,��ci	rן2�b�LD��ȷ�q�ZBЊ�;��Y2��ua�"��F�\A��ՙ�#�l��T@ȅ(��:�j��cb�4`�0�\=\)�$�x\�#N�4��љ���~ܖfb�W�L���{�vQ�Ə<3�9�/��t
��T���p����%V6yخ�>�|Oi蝁}�j`}��|x�����靧5$Z�S�CI��LD_�N�ـg<��j���!��B�c�Xy��feo����%|�`_�]߆߯S:*f��%�~!���-y$ԭ��TH�s\���<�\k-��$�ڛv��i�*pst��Pj>Sgn�b��C,ezD���Ƽt�� S�I�;=z�G�ї7jF"�Oeeqή��ڑz<^���u��5�.۲l0i6(�PʦѮrb���-T��X=���^����7mk!����˭ ��PI=$���u�uI}�s���	 �ڴ-y���[RM0)_�zR]ص���� �A�F٤��/���C��E�Q���º�L{����3���z�����)�v̆�wdn�b)��'�y�Y���H���
m��0�ũs&[i���O������f��w9|�Vg7 W
L��@vK�Մ>S���;=�څ|�K����&���8ب[l=�"����>������y,����Gބ����^�̠�$`�/s��T����v�b��l���[��-�+�mȰ3�$�,�`�@��lM�ݬ�0.9�0DUt���kf(��4~Rz���:xC�AC��kPxq����m���m��@a�'�u�[�l�6��<��to��y�a� ]�T�*�H�%���>˓05r���`����ɇr��m�2�.��hP �6<x(JXΠ�t5#-��T��=2����о����.Oh���F:���Z��W���r�*`|�c�3�Jb�+�G,�w��������0DGrA-1�7���l|Y*!?z���
a�����I��ԞDE+#|�������1�1<�`|Y�C���>4a����%�;�������}�<;���bt;+�u��0ŏ�cPZr��Q�2ln*YB�����ݝ�����-Zg׳�9���b�Żo�n��v��8���n��B�\\ k�#N��Ň4A�	աVٮ'nf�m�����-���BB�c��-�y~���(�#xO�h��-i hS�l�^�5��4Ie��=c^ql�?��
{ �
n��|+8d�r�$�3@����֧���{�C�S^�����k�c^�1�8x�[�M��9/��E�"�+ �B��^��9��*�ԖV�7�2��9�o��B6���?�m�-E|������gx+�VR��a�� #�eoE���8_���ְ�R~����}��3m \,MS���f��oı�Z�Ib�8�oW�l�ն�,լ�˅��K�G�>�}e�S���v��(8�nv���2�観h���զD:�VJ���d�3�ɗo�eR���1��&�bJG��pC�S�)��@	0�A�2�z8~!����J��&�v%��]�~W���i^}�-8���l�e ���ܷ�E�W�����S.݉�t%N^.2�����PHb>�|[��?���;��Rfq�J¿��x"����ӺG�%qbQ=H���������MP���Jhde���&�,���^�x ��nԚtZr�{&�-D�bzZ�����q��']�˿�L���"�~��M�
V�L(�bc����r�	�)M�I����|+������	%+����C���XŖ��KKFq�����Ӣ�EX�w[�P�"+(f�=�����m�ɤ�t���� �,"	X�ë`�5N�;e4�3�V�o��uy�T�y�� �����d2�'Z���Z=�ADs�s�
��o|3ᶠ���yOU�#�Š��J��YV��j�,Jy�*ο����E-9���ǈ7���ZK#�<Agݫ><�8� =>��cq���**dƳi��S�G��a�E��@+6��g�����4:R�z�=� ����"��b��wu��W���;V	��#Sm���q
_����o?6�o�N]�V�=��e=�2�P��Y�����p�/h�|B��2�N4&�f�����)��Ԕ��M}D����wMмk��eF����YJK���U<���n��d}��=,�"�����nD$�ɀk/X�.�]b׬�O�F2=��g���r���쨆wq}�(��:�#�!�c'��}/�YLg.)٥JJ)�o���,y�4��nɪ�	���L�������Nr��``��d���Q�����?�k{�o��D�ve*Q���f}e�}n�uS�����֦����ړ� ���ʣ;��U܆��1#v�aj�d�;��ؖ$o�.��	x�6�U�	b�78G�3���KˢQ� _ e~�t�)�4]6(�����il��?�@�lDM:����e2��#��i�Ӊ�w�mP�A5h"e�̃�&ѱ�O.H��U�Z�2'Uf]���oC�I��<� �����R�Pʍ���6��8$ 5�2%�17��Y�����ת~������6���@��%K!��}���-�� ���(��d��F"�K/��=�0�ȑ�^��8�[�����P�?��C�DzK�7��EM-z�D��FV��s�b�eK�}���Pᾼ�̛\<9�7�&�!������1���0uEF+���͖¾�]�~��q-a�
��T�b��=���Bcȫ�>�~�Z�0Z�q�5B6 )�f#2��sNTr�n��աFL��t�u�S�Lչ�"R��A]�r�7@H�NWw��X�:�>��B�/JT�G.��p�a����R��c������{�]�~<C@�0{�l��	��H.�<�K�	����'D�\_�	q]�S�;<���4h�t�����{3��?������y[E���l���W!��8�s  ��"��ɖc�����@<)r�3H>y���".�D�Ì�p?g�-�"���)}bq�_��-�|e=��m��Ie�	e?u�Ԝ�i?����Y�o�����jNir;��s��8�Z���G��ݕIr�{gNE,�`̏�<��A��΍c�5��&Ds��r��a��9	D�����:Dx����
�*�?%�%�EMx*^{�\/ ��'�����ױ�$_�;x��عF�:U.���� �(p�I<R��t�=y�g�t�߹"�
E��C7)y\и�r�dģ#(����*=���,O�x���Iw[~0a�L^l��O�0>�Q�U���ℓ��S���v�(��!}��!*c���^=f����߼���_R�ڶ���u'U�/��S��1%�H�t5��]S0�I��J��0n��s��^c'C-��ʑ��}����Q_�i;Ъ����X���xâ+��P�%��T�9p���yHfa��ہG ���B�g���,zg��P�H�I�#�DQ��k�	���Ri�g��(�p����7�M^|���b�p
I��bz��\htG������_ڵ�j�S7aI�j��5Z��v���&O��qi�-�LV�K�Ԩ=�/bϠ%�p����G��H8�x�4��ke������@��'oк8#�^��Xy"����1�1�����`���(fV��4�؃��njĚ&��G'�p1G'@��-s�S�KU.\��-{>g�����{�<(h��>tR�mk���j$�x2�u�"Uz����O��'���3�-c��U}�+W��%��,L�*|��XA˓�M�{��:e�sV��ś�ڨA�ߵN��&�k��]L�.Z�Ou��>J�B�D�u,�ĵ��I�Et�ʔtjڎ
��`��f�������8Ws�3�3���@o�Cf��!�w[���v�Io��^���C�7c���ly\�?7�Dn<��0�OJo�<�A�d���?��#�I\T{��g���84Xm�̓j���B�(�F�XIUGH���gW	��� �|8���Kk�7����=N�wx�9k�]��"�{�ȳl���@4w̎�ķzA�_B�a��w�I~<���(֣)U��Ea��f�/}6Q
����߈6��-�������}�}��С$�tWk�m�<}�[O���9���"ꍩM�H9@�B�C�������M�����u��]`�&`~�5 �o��ךD���b��5J&���g"��=b��s	�>gH�cy>�C>��b%��sƜlҐ����6�8go�uvD�%�*�0Q� �[���yb� }��.v�"�#�8��E�wqE�q~�]\�#���4OLX�����J�B\a#�2��x��D���� ����~$�HYh�L�Df�Z(�Y��h=�9ى�M'�|Y� ��8�2���}���V6f�k���b��m��?�Se&��*�Btt-܈�Ž�l�״�p-�`YT6�|6��O����U@۴���e C 3(}yX� ��b�=Lx$��`���)��ݨu�lh�|N"�q�n�T��Lx yC�sn��t,/Y�Y@Ƒj0��_<'bs��!-���KH�?�#��6��p�dn�~����@N8ܾ��dۨ�(O ��(_6�1�W%x�ӳt�%��[����C�����&�ez+�>�������zn�'��g�!�sO�(�'@T���&��f�IFD�{=N��e/��d��)d���-[z�J�%l���_�&����3��kT��0q
�O��&ѝ�|��A�h?,�<�d,5��8k' T��V� �3ϫT���! ��Y���,���r�c��-6�/<�i���CL��i =��j��wf�m��;q�~'�;�G�7�+ZkE�\ 	z��1#?ߣ��c����%i�a(��/5j�˜_��Y
!VE�O%F�ys���*zEҀ�ˠt/��1����xNI�A�ӹ�M�4h���'[k���}ޭ�J.K?"����ki��4��5|[C�{]��g�@˛�H
K�u�~P���$'_[ZU�x������T�sN�<w����u��ػMh&�Θ��!?�A�&m�vI���R��	Y�atœ�lc��CÛ�І��տ��"���_�h��b@Z~pr�|�+�k�N�
x�h�i~;R�|䂙�p�+��[���O�)ׅ�m9�Q��1��G���7:��b1�G	�Ht�����a��H`�Z�0�:�1���q��Ym�����l�Z{̂�3*�"��Kv)ψ�Vc�W·C>�CW�+����Ѧ,)��3<��96D��OA��P�-r��&�_�3j�=a�Շ{t�i�'Ֆt���4����p�-��q��E(t]�!b�4&D�0��@K&Z����8��xf����M�����6@�D]�j�$y5`%������n�9a_M	̣>���b^J�v��C_�K�J� �=s���{Z���:9�{Tc�׾g�AF>2�m�A�ܖ�-as��aIu�*�RV���UQ�o����0D_x��]���vB]�釞[��Ԁ_O9�X�ȓ2p�D�����#�p�ƪ�I�?g_�8��g���0y���kj��b�x�l
Y�?�Ic����Rm`���$.͋ʹ��s٥vFe��>/
�D��[h���W9*�q4�-��F�{/"���<>ϲ�x�2�;�J�s�fd]��x<�6�6�����tU��� @!���i�D0�t���d�<hُ�J�O�¡���q_o�AKpҲ/�-9蛊�1<t�E;�IJ�x�!��X�3��cQ�A� *s)��W��F�t�u�|��7|#�2W���ж
X#�G�g��<��<�1vn��3*��������I�u
[�g���.���-��Uw�OJ�)�w��`�z��[���^=._��W�;ݚ�'��������v�;V�8�K��>��t��jƮ#K3#��3�Bj��Ae��3��Z��W5�~q}��"e�I�������Ѳ�Lϓ��k�Ov���Ai�EG��n3��uk0��@��s�ƚ4�f`ҍ>�s�W��Q�p����Q9���h6yJO�YjHj�l���C�ĸ�,l�/:}�.H�'�ֻb�]V�����U܃+�K��g�0��]��КJ# �3�O����\νD���J�.��/����ߓ���8ن�ۙ�6jP��b��F`�u���@ad�-�J�Շ��J�8�V�E�Z}�l{�cK��cn��<�ܔ�oE;�8uiJ�v�QQ�Kv�Їv�;;ۺ0�|ԩU1њ�L2�R�������1ӵ��r�e��!꨼�K�1?��}�͝���j�p��5������62�+v��4��6>£�+�?�'K<;�KO�u�lI��ܳY>�� ��^\��=4NY��9����퍈���s�")�a�x��NFI���E����kL�h�g�MWZm��R��PJV��5�c����43��ĕ,o����+��6Shz�MS��~�nN��a���6�����5s�'�����]�T��I��}M	Ǜ��1Tk���
g��Cl��)�s�/es��dTⱚ�A:��N Y�IN����rKa�$K�Ul�Ԫ��jrޖE���`�2�bsD5M��B tAg�_
�c��͢���hs�1��Z����@��P$���QO ��6���o�dq_	C��EҨ?��$B�!�B����M�����y���g��v+�L���U�A_J�z��T�^E�jT��t*z:�K_�N�������0��p�����i�r��oƧ� �gUIځ��P���h�{����K}����Ȫ�n��a�Y]����!�r���vQ�
`R&�{領Se�]�h�v��x�)Ra*+�kKI����Y8�aH)|3
�of����3o|M�ףuu��iNY��A`���N�9�$`ܿ�Fm R���W~kt���S��[>]i3�o���n�4w<�@	-�����\�:sUqAhȘ�h�n�1<OwnɎ���T"[�D}���}2�<Ě�s��a�e���>��N۶	P�����7�%~l2�A���r�?�d���`���K~��V�A�$��i�����3<�G��ng���|R��Ά1f�Ѻ�8/z�28�#�H�S��Z���M�:4z�%�~�wt�IM`��#�/����lH�d�v�@���c}�>q�du��G���s��+q1w.��
P�W�X`4U{���_�
{N�6U��D�;n��v�楃Ƶu�*��^�*W6<�o*-/���w}���2��@���eꤱ&�\�����~o9h���.��P}����ښ2�����Ԥ������G\r��5�ҶF�3���,��9��$����D�)��7E#�Z��ђ�a�@�Ā!*˹-@9��IZ�7�ނ�{%nrY}��B��v�J�-�-mI�-���u���h��	�km�����ia}����@�V�4
�?���d����s*��m�y�/���Bʳ������V�#H�p0u�h>6����x��[j���ޔ���ڸ_��ax����
����� ���Ap�o7e]Ǿ7T�2 ��e���3��7_ި�ހ�=d�6�ȸ��O<�u7Ώ�§ĭ�ꗿyӀ��@�ps�ٱ��f�Q�����d�&k�ԹA�;H��@��Y�9�t�A�r<�}ON���+�G(�,����;!+eD$��xeHq�����&��\,�'�T��F�ٜ���%ʀq�E[|v�-7\�_�Lڑ��:�y�e:��Df��biE��OT�2�:埚8#,%��(�S&��v��te|R�i���D� ��Yĺ�
u������%�_�S�m6%�k����R�нs��$i�/�W�w�| 8z ��qͼQt���=�3��h����\ؙ��M����
�5G8S�<yfN�8Lx�H2g���nT����� ����h@�!0,�1d}~��
E0����0��V�hg3x��������+u2Ϳ�k����$𰮱0	�J�ei2�����}�CFS+���x
�����uĬM��4�4S<�x�E�����F�mx���N���e��|��V��紏�C�O�m4��3�æ&�S]�0�nF���Y_�_�g�A݅�zL���a�.����296�9�ğ r����.�*�E<6&�R��lt�H�k,���+0�D������;na�>�&�3�B�̒o��$�s,�ҵjV)0O�V�5�<Y�3���o��~"s���d8��� .��$:m;�T<��I�VWڭ������z��2��d�1�H���z?ru���>�L�ᒬ�c�\��sޅ�/2<�GOt�h����*����X;wh���V	���'��I ���g�D �j�֍R~�ء�=�su�_����d�?\r��V�s`��\�������;�P��T5�x�-�(���'UT�e<F��O�`Q#~���7rs�RG �ShIb�Ok���'���`\�<y��V=>[ܑ�n�|�JL�T�;1�����a5�g�FZ'M�R�d��L�*tʃ�Ltd�9X���Upֻ�K��z��k�m��Z��R-?�]��jPF6��R�?�$xAi�Ơ_3�>v[\�<܏�(wv�1�ı����s��N�w��|El�����zfm�fJ�����h�\`��?ҧ:B����� ��S���R�E=�p ]=�{N_�����Y������"C5�U�9R�����}�VbX���f4�� ��L�>�1{(���T�84 ���ڪp��{�5�����ݷ%�׌�ad��<&o�a�����Oͩ��s�]��D��#s�[]��	�Am���֌�lh�zw"h�p[S'��{v�g�`�۞�l8t�LyLMC��YR��~u�>��z��3Κ�*6=���_fpw��I���8y��L��$E0�y6(lz�����v���^�X�kݿV"���Z�GpX���Ӕ�w-I3�z%J0�w����c��	�&d����᝟AUZP� �s���& V��%���3!�TRu�Jx9}��B�p�5	0���#���N��e��L�F�F��q�}Qa��9a��~ٲA�҅�_v��~�]&8�0i�\2؉�w��^-������N϶�\V��Xe��/`�[����X�x�(.�H�x!P��a^;(:%+�/o6q]v3m�і�WIȢ�x�\r�b���"��r'N ���85�ӕ�v,h�Sk�|��P�j���N��;啊
��s �V�m<�w��7���K*<�]1z0���j)�t:��n���}I��ط,��<]L��ki|ӂ�Y/�B���_u�j��kဣ��� ��NvH��>f�ɭ�&��h���?������C��2�)㩳���8�&-�޷H����%��Wwp���j|������OˍV40�]�ޟ�O���_n-R����O���v� C8�����Q�%��ܸ�6��t,3]�l�!��k�Js�!���'���}�@��.Dn"f2w�5ͯ��ZU���?c�Նu�9����!�i|-"]�n˦'c�ع�loFQj��b@3�ũ����Bca��[\U��:S'n����we?*�~�-�{��H�>�1JhIR1b��@H��8>bK�s�I��vfF�{���l�2��m�;�V[�U5��i���G7UÜ {��z��Ͻ�[�~���.�����\`>e�pc�*�0�����FoA�K��e��[�t���X��L \��s��ҋ�B��"i�M���dF�M;K�M�*@09�q�5(r�wf�]��ъu�����+:~�5"�^���W�F�޹���!��nH��K�����H���l�'���_�� ��	G���Q�X�� V��Zq�����+�q�с���U��ʦE��YW�yBg�����ŰkP���8�5a�Ɩ�d���y���B8=���������M�(*�X���l�v��OP~�WA���j�������e���%ѬFF�(=�y��='zJ,Y��g��~s�P�F��!ސRL*���4�0�$*�wV"Om�n�i~k_�B-t��@��HZ/��$F���!+��X�D�{���g���Md��I�M����4*���Fz��
�B�������7�Z�i�@��ە� V4zz^�]��ӽ�DQ�{Z%��#D�@i���>���(��	�~F������v�!�����^-#E`d�t�pS�0�J�َ�"���IV=�w��w<�yD���>���2y&4� ��i��	��ȗ<O�%MD<� ��g��4f�i(�r�'�Uw�ݭb��4s�����g�2<,�5��?�1���T�ی��CKn6x�b��vMv��Ӈ��K��'�Kz,l�߬4��lՖR�f�{g�����f�H��}����c'��V����q}e��z���m,_���Q۫��
�0����Yض֍=���2��sP>�����M�rU+6���C�_���1a�њs�=�u���sa6,�T7o��3ȸ�A��2m��N�לqjꞟ�;�u���}2�L���j*��pF�)��G��2�q�K��G���/���K�����Պ�e�i�U�'K*uN�DOg��H� ��Z�H���@r�ݱ��f�R�>�Q�2d��uX��9͡��d��H���׵��/G����sɇ�(�� �\o�Uf3�3�V�[��óV�3��N�]#�FzgP$�tR���5R�:���<o�>�ϋS�8�&]!�Q�F�q9h�x�
P�V������ S�)ԃ=��يtǙbj
����:iC����7�p��4㒎�@��"�'8���_b���K���ǵ,)���C�4��Gz���;��������^2V�1@��C���;y��;��t�b?吥'kҭ�|2�^6���1���B��mv4�n�y�'�q�y#c��T���W#����?X�ĺC���̼_�d����?��~��p�2�.����,/Ru-o�ϔ�x�W䡝�>�F�OL�%.�23=��T;	ɇV�hD`�S�����) �������T�G$�����W� |j�_̲������+�a�k��ĥ^��pK�B�A�q��x!�"�wf�h�M�g+i�A9�$�A��.��_���$Z�y�����'���uٖ'���uh�5��s�&���΃��ֽ�
��I^d�}͸�Ef���0w���a����ֱ�}�zZ�e�i��ow���5`9�5㲢`=�·\�O|8B��w�u��]\����n\A���j�������diR	�0�����{�#6��"��K32f�e��I䍱SP��[,�~�K'�d�-Z_��S��r��|DD�BӨQ��uD:�7
zp%5�DW���y"ve1J�#0���C���/�{<B��Ѩ��k�Z���eoR�˯�5�^��]�-	�5���� �g��xr�ش狲�Q�
�lR���xM`�0i	�_i ��E�#"W������0��I�=� [����	h�a]����xa��_Mp�S�O+<��G�9D�꯱�����o��T��!��+��So�y�� �7p�b2������	ƍ��M��[���g �$G ��<�`�{��BϹ���tZv$D-�X��N�,V/���0d�}v΅��#� �Ƨ�����EEL��c�W��?q��G�1���a_�d5�|sV����J�<&(jm�X��J�\�C����N�+�'���0����>Q�ă�ĭn)�Ǒ؈�l�!�a��dS["ӄiׄ8=b�Yl^���3�!鯈r�6͂��S�W*	"��Q��FrQP�3/U��ʁ�`|F3L��e0��������g	��[���=���BZ��0��e^�����Ej�M�t:�r3i��������L��.��z����u�M�;W5l�U<����T����΋|�e8���2Ae����;)�uA$/��Z���p�?b�~^٨fM{�f��Y~�j�s5�`�7!�6�v+�$�Wɰ��YY�1�:�'I�s���ܮ��o����c���D6���4�RN�-���qZ� ��$�vO��M��zg,�rd��<����l�ShL�t,�(BMG�Rܺ�@fL��뎬O���Ef�O�&_�~��{�vw�)�R�/x��z�0߽�H�m`1��^���wF�#JuvՓ�W���H�
D�D�D�e�d���ɂ
ź��1���s$F��OQ���lO�#��
���"�6��*���g�����_�ugw���#A��e�J�l�hN�~φ��������;<s�A$O~���~C覨f"���7(]Uj&o�B[1���&�V��ҳ�o
�f�1���8�$��!0����S똋���9
�S�J�<�C��C��+$U��n�:��o�Q�T�\#2+?%�l��7�"Ăjz� ��ʜ�������" ���o����gg��F�?���Fe?p�.j��ے��ƹ�ih�a�S��!%��@ѧ����͒\�g�Uz�*�[vwe��$�D�.�66@{���^��x����vJo~�ʣ$�3�QB�8XE��_��Bd<�����2]�=K)E�K�]��.Z0��:C���t`�o�G�s.{fB���+��u|.aQ���&9�}����--(�ң"S�&fRʩ70�K*�һ�r��6��ձ-�ѝQ��$#��:�0�@3�GQK1i��E>[0ҧd'�:����%�/q�c~<�s��s�����F��h���}ܑ��9R��5�Ƨ}���|=��|�f~4ݡ%����Ւ��A��;;m��3��Wj�`Mzdc��,Z��	̨ E�����1>�tF��2�k�Y岚�X�p�Y+!~EO�Ȁ��S~^4K9#��(�J*�V�|1��&�2O�7"ۈa��o��t �
�� "=H#_�	�ɺ�5��Pa�r@��5z���9)~[�X���}s��r[�iz4?�ö^���Zu��������c���L��c����d@�q�J~����$'��A_���m���i��>Yh�2�5#��G�B�#�Z�4r�D���Q]��M�@gsT�����k��I�b�� 96BŃ��G(���W��?$Ip�P�y%J�7���+�P�y���/�p 6\Fl6I7��T�E��Kq��SL�V@UiV�4�U	��s�pܤlLvْ�*�}�{�. ��P�靪�)@�Z��^�R5��.V��{Ӳ�P���8��n@9t���w��L�h��Q��3h @1)+x�x�ªb�n�(/��F��!���脀��~�s��xˢ�"b �E���l�B\6/���s�3�Ǡ+�OX��JF祟��i�Rh��ŗ :?��F����2�gf�f�В�|�����8@��ۻD$�M���].���A/D+�=�.6̀WV�^8{�-N�`�䜐�c���_^p�^���?/���LO���)0��ҥ'�4����R�o�刱ЁUq����̓ҫ|�A��s��!��p8��]�/��;}��(��"���oMB�*ehAߜ����8�w\�r����:�V%�h������F������`K��<�"�m�2b:{�!Q�O;E��$]�j���C�U1,��J9�*#�/'���oj����P�܎��FV�F~�[ӳz嵅�P�"�vO��,��������5U0�ȼ�m��Sl����խ�?/P	[��@Oq+��_���'�.�e�eG�����9���r���a���)�GNu|B����L�M#���z@|�f�m=ĝ����Ed�����K"J���ƒ��
L}���;����D�I����Ax�B�}x)/���j舍3w��~�AV'�,�Y������~��91���a[�4�`�>z�o]ig[�{0���ȵ�Wz=��gI a�jy'ݛߥ����OcR^��`Q��;��c ۑy�1X'�����4o�AE,LK����ޘV#�G�J&!�	9n�I1����$��>�D��=
������~��]t��W/�r��ox�&��ח�\�B�ZINq2Qi_uׯ;�ȝ��6��s(Z}ԁ�
��y��1І�7����!݅�D"�7�� L���M�G���%�9g���QOp�r�}�'|�s�7#k��B����aP���u1�h�'Á�(�t����X�h�9B���VP�e����qoWӈ�9������"�tV�BQ����������s)f]Z?�!O��	S��h.v��A��C��� �����P�#����(�2��2>ޕw$ֻPf�&/틴��֧0�꼴(e�2L���~z&�Q<�m(�C���Y�@�U��mU�D�TI<<�X=9f��ɌC�Z'��L��<jm@$�J������:k�'���z?�w-m>lq��>R_�S��<F��V; Zs�M|k]kѠ�!�Lo�
��b����ض�δ�,_5_�l&~�sL�N�n�]��6R�4a���Q�zfF�����{�Ɂ�3�O ���]-e�Y���:�&�pap�7������m�7
.-	
Z�����?Mֻ�����Y�����݀w���s������)��^��̫`���0��n�G�M*�"d*���ԣ��h�
�u�}m��Z�n�(њa���ܷ-xJCƙK�[v�XƆ��.�M��`���of݄�Ltyv��h��� 8z	�W=��h,��-�{�c�D�ߓ�MP|�?'�O+�:#E1����ؘR�t��ɛÎ��x!)�{� (�?;
a�n��.ݎt�5���W����ǥ�1��t#����S��?H����s9�����8�\B�{��_5�����6�.��n��̶ŜM��J#J�SU}�u�J�g��:37pT�L4�1��M��N���vp���°ET�yة-M�L�Ӥ	���:�#���)��w�-�y�`�P��R�D��{E_�����\�ܙ���j9�ʵ\�$ۍ{��|���kh�����MTr향�n�G��t�t���
s�U��<<�<q�-vr�ΰ��a��|��x�����E��R�f����?���u�Ӕ�}���Ll��7�L�ܵ��a%�~��CR\�_�(��#t�� ��[i@d&4�~N�0>΍�TDV��8 Ɓ�4AK��Zx�� �vX���b?6�9/�`�v���k�!���A��湔����e�ǀ��C.-��q	�$8(ؓ[�S��� Q�*�qͮ��1-0B��{Q�o��]+r%���d�E��I�x�ZS:\,�D6����>8�ڍ2�Z�6Oa,ޚ�|/��t�ӜY	�!4vU�
�Y�dO�r>�w���Yw?�����	'
��8�|� �Z6ށ#P�z������Z�5�׏%R��vk��7�
��K�1��No�_f` Rˍ�q�3j��h����lє�ћZ�X��=���1�or��y'����QO������a�Ɉ(�wJ�P��XvM��E��&h�P���C��ۗ�0��A��ً[R��o`E�<p��:$�d��Q"D�4/�{Jq�:���J(���p����#���#��=�����kR��/��S�U�Je~`x}�`do���_�����Bv���L����ꈖ�ė��ߌ9�}K��\��;j��nAJ���b3���*4T2�/�E��H�G��}]�k�]7V��7��DT@���jmřj����(�}�i@׺@�l��"��T`h����6&}L�*/��f>�eMڻ������E��#rL���7���� �G*�\-/�)����W�JH�� }���*>�v��W�[S���xgK	y��i3�X�K0J�� �
B��n�|j��%�z���2-a���VC�P���yڝOjo��7ީ8:�u����"4-���]m���3���\���}�eW�	�ЩX��4%�nj�P>��<J����탪Z<^�-��Qe��$����/��Be^y�`���%�nXv����t��k���`�z������D�h9d[�� l�N���J��iY�t]��P�Ĝ���Js>�M��s�N�d|&'l>�5v����f�┇�k~&�}ba��!C��T�����*���V��{���푝��@��٠I��ʕo��\�����w@��� ���:!��݌�G����Fͳ!I�.W� ڎ`���9�M����&���(����v�ՁC�ْ�\�E]O�3��oMȋϙo�����x��l�M宇��d
���^'-��h���� �*��Ɇ>�t���E������S�8<>�LW��!�9��|�yH \��qJLخ�?�hT�=��zWa�57F��En�Qݔm����v�E
�Z�]M7VL��܈Pu0|��a��E7�Ez/�K7��.�"�Y� ٭��6��!�wM�3W������e�2ԛj���FK���+^��lX�?��f[.ȳ4�.=7}:Hg_�M�? "bc�E��x�M{�e�ѨK�	���Ј�̑byap�!�h.V�p���%���8�s5���������Q��5)殛�r��U�"#?�+����L�5Q�e�<w�rO�I�~b�+��	�"���$	�>g��8$�\�:�:(�i_X2��6Q8jɶe;����Y
)�k�N��̪�+g�(e{�F�� 2iSrjJ����E��h�e���[��{�;��3@�{&�W�k��y���m�Ya-S��c�V��B?"��$�l�W�B�����oy���i�	�m�Z��8�qA)�D�f�
�ȱ�o��3�C��G���ZFh��u�S��#I��htV�'���ǇԪ�v^�?
��p�3�Q���o�s�\��ll:��� �~�M�B0��"��ۚ��e��3�� �6�dgW�m	��ά�l��غ�q�ًH+��FIqT�
C3w��,5���!��$�VܘE%�����O�\K��o��*_,LkH�蔠\���W��v���{v��"����e)+�t+A��!@�z��'�a�N��@Qh�g,�IY�{;;�d�����1a���p�)c��y�ٿ	��~g����H;���E�e�H�&y�#���O�/��Cb&:,�",砌���d|E��Ny*42MM�t��M$�Jo��E5�~�J}){%��8b�3���־k��;I}�����A,m�#�`�s����Ĳ����X�{.gXH}���6S(�
� �BF���8ɹ����P��$��Xb�K�/v���P����*'��Jɣ��?�g���_0��}�,���2�P8���(��)��'���zCTu���'~tN���֡'G�kCqqE�*����>4����� u���uZ�ړ� ��<�|ɼ�w����� ��@z(�g����`&|Ro��ĹM�Ǒn6������u���WU,p2}ِ�⋝��6X�C��?�� ?;K�#��۞E�f_�9�!�;��$.�5���%e����OaN���aJY���+[)݅��%k�*AI��Ъ�ےgět�	iޚ�j`�k�ω������<�����[��x##�ǭ�+���?�����D�@�2ą�.��x���n�6v�x�no����Ñ�{�P������ w�Ӭ->W�[��\j��פY�K.m�
&�̅�]�
S��b���(��|����䟿x�GB2i3�|?c^Z��9G����!~H�m����U{���s�[�Y^-ױr�s"��cv�YNA�)y,A��ȷ� O����a�yL����1G�y+� ��"�4S�D~�Hy��m�C�����O��Uèq�.m�B_�XB
gN x� �^�/�-�%B��l�;�����W%�b��?�v�t*����[ܘ�	if�zn�l���0U���x},r٩y=��U�AQ�/����
��#���M�7��h$��rO�۩��D����)���g�U��B��4ZUbE'��sK��_6��F�(տ��Rǲ�ix�lD���h ��BƧt�|�����R�'�qԀ��(T����S$�@K��`~-(��"3�:R�=�@�������
W�T�,Y#4��G��H,�@�[��۝��x������v�ʰׅc�8�f����y�˅&G}{I�E�Oɓ�'�����)�C:��eJB�<���V_�K1�u���b������9��,�&d�\*�mT�:��X�ꗯ�m���y��v�/��*3<�ft�d�<�i\���c��CJ���+�y�8�S�p�?�$0�"��
���Uκ-�5�iX��pd���p=p���PRJ�R����n)����f���r�>8�ݼB'�;��E���DEP0���<�#+� w���Ic&>�]`���)p��4C���˕�M8X�0�)k��!�&���?7d�VO��¤P���c!S�U��3��X�&,"��Z�2����df�I)[��{K�l��&�ڳ��rS����l�ßL}s��T����(}2��;1;����J��6��\�&�����R�������G�z�m��BG��/B�T�F��0q�����j5\����.�Ӥ� ��N.)�Z� ���H�Ə�h���hh�
��u�I
�f3��ClΩ�rFd]=v�����S�y��X���kv���4Bm��1W�^A��h�G��Z���x������B&����\o-�
����o���b����$��m���zS'�]��Ϧ�m�d)t,�@�C�ϖF��=�J�Ł�ߪ�@���	a)N:��|Z6�Ek���:SUݞ��v��{�(!���p��7�g�66�T3���OB ���!0��=?�!*���/�噔���p�;��ړ���� �W�(\r�p\t�GS�N*�AV�2�A��	�fb�7�ZaK��%9����py֛ Y�~�BU�$�OHhC.^�g$��zu��R����x0��M���Yy0CF�����T�F���o�!=ףcm�!/���h�s����U^�r�
.�oΆ.��%o¶�i��9tȻ뤳҈�o�mJJY֓c"��,t).���\:�Y�.x�G.��3|���^=@����J��.�K����{Ws���;�J���60���/��ts,��)50�u��F�^�V���)��%=�=KS���B�����M��Gh*�c�G��������w�������������\b`\��^��q��A�!�4���I��"�H�m��$����Ck�5a�ĉޮ�,�'�pbe�j�(�xC'������1��Ԕ��x�.��%�{�D�Ξ���
�`�I�"�qx��b��S뻫����8ծ���#_��#�r��]
���?*��c?��4[���k��Z1gV��m��ۆ(+K�Z�t�Ԕ�B�uc�2c��HO����B�z��u��	���0©*���dF����B&^�<�w��xT�5G3���wSX�%f�7.�yt�Bh>�U=��Q��C#���[*f7�pp#"����}�7�{�Z�fꭳ�I�O����
���BI78I¨+K�����Z�.��7���c,�m���0�'��پ=0>rL!��f~�x��KU#��bR>t�/�'Ǻ�t����W�L�}RJ}��g]8�6l1~����o��q��W�U���$[��5DZ���S�������͐����`�2@Z�~�v���l���"�W�*D]�I���bǊ�����篯O5� (��V `����t�G�o�&U�p�=��Dv@�>^��8�3o.�|���6R�a�"����l����cJA���]��,R���Ju~�6�u�ׁ�N:7�*uՏK�����>;Ȍ$�@�O2��l�`�x�$	���w���A��?�)�Y�,Pa+/���t,q/r��<���NRg��տp�u�z����Mc#6ǰ*m��_�չ�R$�+ᦌ�쳏|g�#_�B]�`hm�k�yJy��8ށe��JH]2u4L�E���	P���Ou�U��� XV3�_�m��.�"�8@�y��@]΍$;Qp�A�Q���#�6E�bIX�Gێ��`;�YrOHЬ8����a6]31�*B�0z�H�����НI��}!��=�O�wЩк�E�EC�uVW�G�M�H4	�=F�P~8���<���>A�:����`��e��J��dl������H<髷�1c3��ѫ�k#�#�m緀�Vm�&�F�%/�x�J0���m�t���E���+��6�U���+8�3p@,},����l�H��B�+����I�.��h:^ijS(�
�g�U��}y�/#gp�t�#��AF���Z�i��pI���QU�Lv+�!�A0�hu�C¶g#_8,���B�o���ewc>i�[�8w33TpIPE����L�o�;�m��c��32�]��3�>s�j�;N��TZ�o�K�2~��$��ya��+����r��V�u���޿V�Ǧ�p�xY{������â-V:$SW�+��>�ix-�-Ƭi������l
��I�&#�^"M���&�c���k>�AF���b"^�Ԉ����qL�;/d/�,��Z�Wq�W����G��3�.�;b��mM
)���/\ ��+/����*-5]���d����E�^#k�r�t�G��&�������Q����$�l�B�i鄡���"��p�h{P�<g /`u��E_I|S�-Ɠ��D���[��\Ͻ�K�W?Ɗ���$NG�w*H{�25�V#�X�^uv��?j�_�}�X����Y�-��0��~�}�j�\i-���~���
����"�ћ�����v5i�tIA^���H-p� `��f�< �}��ԗ+���$�8�y:]"@(��d*�wv|�۳kܠ�1����?<��z��D���SS;�������s�m��Y�nŎ�J^�2��if�Aai��}��#R6�T:>�DI�t�@�k	��e$!
�[�^�\�%`���`�B���ef���S�h�c+��|6�+�Z$\f���A�`=���~�jWfp0;>ZS��6��`�;K��$��ýo��n%����m��ξӫ}��fx�Q�p�t/Z�@��`��� �gGy����z(�Eǟ#�~2Óq�f���#ԡW:*�"���4(�Tx��ظ�}��l��.{B��%��݀!Z����`7��"�	�o5�1G1����˵sc_Ģ����Q�AĔ��I�O�!��G �)4%0Yd���� y������[��#�4�m�y&i����_��jͩ�bK"�(��e���K\W`�$�wy���Ơ�A*7��Mx���=�Ff�yxTn��j���-�$�\V��.��A�T��ݶ-����e�A(�`���\tQr��&� í�Ym��7�t��������H�@���a�$����`�n��P@P��.N�ֳΏ��Zcp�,��+Ik���YTR�6��Cx.��QeME>&�l�uP����()}�XCR�ߕ��*?\���\	`�e���_�bq� :��_�˧�Q"�k�*�E�2-w��':"l�`����& @aT"̯-zw�FHg�ؠO�ǋ2#d��g���zi�J�}�U˜R���p<�YA�W�X�{H�Jp�%�a�짝*���<�0���2l�B�ʭXΏ�5{�PR��F��ܘS�:�M��|�7ȧ�ҥbT�b�|��4�DI�%�O��H��F;���tJ�~y�Ů�P�O��R��IT�?�U����!,�]�����b
L��'�7�yK��nnn��1:ߥ����;:f�.<i��R�~�h؄�^
�X�y��Z�����E0s3n�8Oo�����vC�)@�1
��d����l�2�����D~�iu��!���������Td�{:-��yu�q;����fEM�Q'7����[ �`�ɢ�'������7�ѡMg	ɥ�T��U��x�@�����ke�X7��rJ!uë%N��;t��B������-�'zD�ֶ�_�	�8��������'��wt��4�
 ������`̝
o���'}�CP���A�3�Q���]S��S�m�'ֿK�?S.��=�|9�2��G_�Q�]y�3�{�fX�FSS�uI�=m�In�o��8@��U���a7�����i]*3	_��-V��e��һ<���0�ܣ��ݰ!d��"c��Ģ������ո�	�G����.Φ�� ���P�ܝ��R^�����⣴�i=���@*�+xAI����*����G����&&�<t��*�?�6��}Օ��G�	���XIC�C~��TQNf�[��U���*T�O2+L��0�,D��ަbGgo�������DM�f���e��s�	F�_��wR$�(]�&�*�y=y�������i,W4��G�_�{�0%b�/�4b۟Wǻ�����1�er���p�L�h����|�[��U㐃{�=MW,{��)�s�]�!W�+��ʎxC
uU���7�+K�8�B^�-4ǿҲ�����퐇%톦=� �=������0֯7�2������I��\@�mz�����5��B����G��&r`���8�BT���q�)8��U��/��)�͛�
/��W�3�+̓��R����)\	@�h�$�2茱�Ж�Ei��u�r��v��t�..
��ܼ1�CZ��d,0��-��]�-#M�Hv��#���48�GJ�Н�'$V?g"q���ɭ����Ț*e�-S=.������_���e۷ܬ���ǚ��Z���/��qYJ��EEX�T���8���p�Sy�`h4��	�[�}a���/--q������P]�e�=��8��xG�FoDp_�}o��*K������2ft셧�*MQ�Jo�<as�ah;��\�6���IWF'.A�BH�yP�|Ü��ds/�����4K�oCʡd�� ��>���a�7�OzW�"��蓓5{C�n�,o�"���
���g<�9��((|M#��#h��+w��3$;(�����(��994��26$�z�>�N$�r��8ę�m-Jeke`b4j�����#�D�f��dv�@3=?K$�Y��h�� ���z��T��|��z���D�c&��uԌب�ߥ�]i,^t7�)� E��f�����5�Ͽ-@?/���H�/����m�~���n��°�iWQ?6���-�U�K�iD3a��5��Z�Y7N���D#C����H�X�lP�[5,����O^o~͎[]�JV�HZ��ݢ��z��b�l1��O���G��������Uʳ���S�����2H\��U�
���-�
�a�1̀������ "�syy��$�#8�]���G��Z��.�[�\_w�Zk�K��9QPL4k��Yr��;u'{�B�"݌��a�w�����
�jc����"���C�h� �Q� ��oT��s��F�Km �����CDD�%
�k�o(|���ֲ�'��s�Q.]x#����Q\�#�U�Tf���`ؐZ��""�����#�?_6\EM~������"P��NS�<�/��F��޳z��9*�T@D9u�S�O��5��� �s���Ԃ;#p�q��p�4��t��YPA3
?h��k��d*!��k�'���,���:v�t-��BpH�ɩ�j�[KL�n�B��_�'�����{� [�ߩ��3��ؼjAU�
�b��qOf&�����\Ki�V��������U���]4N�A5|S*�A�ѱ��ͽ����J\��j?B�	��8������TLɱ4�n��9���6Y���*UV$|g���O����I]�DE�n)O�ן	u��=��������tc�"��_�;�W�|��
|O��'d\q�	ID���Ĭ��5�J�:�����&�Zo�P.�R�I>�jK*^�H�֜�5r~� �� ��3A�{���1�O,��`M�sFX鈻l�IϷ����M5/\�oU�,�UU]R蟓��%W<���3�{��i�0#1��Q�ެ�xl(0K�(�D R��O���x��;��l�� P}Q��4k<9p��PH~!Q�%��M�w�;H�����e��R�^��j�%w'����92�4�|�ś�|�}����6�,��u�����@�碇*�LSD"Y�|0��I�̯��?N�RM�hW��Y��U�����'&DU��[�3��`�<���dsu:o��n�}�B/����������3�Ѵ�y�� ���SP��Z��n����]����^:S���Z�u����AVK�d�ٸE�B3����Ø�1H���� �B��=���~��*�c�e�i�c�҃��;ÿ��8�%[���g�?�m��� b�5��R���ñ����q���(8���ᢷ�	<�mT�g;̔H򧚩��8��a�ӀH��J;��� ���;ş����]K�S��������SX9��]J��#̏[&��0��q���G#�Y ����]X��;][�_����S���v���[{A:m��Дy�j�;Ȝ��cZu�,��I��:O��.��B�����dޜ����\���Z,�U[��&VTj����r:�k�u椐��ot�a��\���`�h}��$L=�AV�yg�-�ᘿ��y��!;�-(\��`K���"wL � }=�B��8�\��3"h��[�����3^o�Qa�t�Sͤ0�r�P���+J�ɘ������v�C��M2X����7K��Cǁn����lNh;�T=�9��Á��Լ�V�P�B�W�+��*�l:X&S��q�"���*Y;�_��zNH9k�o�Ur�gZ,C�g#���F0.�i'C�=B��6<�����l�x>�)5������!@r��&DL;��ݚ����e��*��u0��g���ɍ>6d���m��S�h�BCJ��Dq�X�`�:���%G�ѫ�Vg˕u�_�\u��g
�>L$6�Z���K��z$L��H������i�m��YW�xb��_je�6߀�����Z��G��(���	�/U�cFԒ)��g�t��~j�G�z����"�c�bO��>����Şk��M�h���uNf#�]�j��C�%�D�wX���\ȿ�[�{	��+|�Z`��dM�d��6'�_#`Uei�-'���|�Z���cT\�E�L� 15^L����&=�����������J�k��z����uO���GR����QǶ�t��O�b��nw>��������d�e���@d`�&y��&�� J���lɽ���MwZ��
e��R��.|��=�$�_�U�|���H07�X}'��uT�NMB$#�:8�l	gɃp���]�r��2�R����%�g#d#3F溏[A���s�)�%W�k�J}���D�W=��v��|���n0W�'�댲\���������R�*f�?*���ׇ����v���vo���W�j�451�(�sˈ8�~���(QںS�9�TAӢ�װv�n���A�]��Qx��ڡ,�B�O�8�y�	t} 0py"�*7�6�s�a

G���j�͗paE.>����o6���n���D^�B���a
ܱ楅% S�l�Uor�����`�6`��o{k@j�m�1/G=�K^=�T	tlS���eX�lAA�V%d�,n��]�*�"�^�H5��=��yuޔ���W�.-���)@`��Cz�� �_]�)d��2�f��������͐�[�o�H	��|����E˱p
mAO8���JĪ�v�΃{�b-��6i ���z�g��i�v�"�;�SY�,$�o��Z�-�us5�rep���ܒJ���WA���è�~��ǔHU��R������{)Y��kv!>��������.���p���S�H��z�tMʎ8�M6��_�8�2�O��x�j�a�v/����cP�^�����j��g�U_�%E��O���Y� }c��l-�Nol���t��-��wEhV��������@���S�@<L�N�%p ZX�Y%�썬eƁ��y\���b��y�(.+���!*w7��Qǔ�N_�sݘ.�M:qW�͆�P`*)�J1�8mr���p�O$�ʘ�W��d�#�/�&��q�0�Urg���@�'�k$u��Ф�'�H?/��ݙ�E�Č����X�딢���S�#�n)p?H�q��>K���@�Nr��*��KW%���3ϲ�k5�z�sc��F�1Nqk�c��/��E�K��>���ek�/v��dM�¦	�ȕv����ǪR` ��(�L�ǿ��}�k���?��O�����.�&�`X}�}j����ÓǗa���?��7`ٟ
۟*S�ȗA?ퟭ;�+�/P�@�N���e"�U��P�QRIj�N�/Wk;oItw�`���`5M�+�"��ak�]��(�dۻqHs����Eɀ�s��������?�T�7��WG]X�"vf��F���3�P����3>�����O�Ӱ1=)GL��	9��b��P}��N��
�ڇ���p#��u��R�d9�>�^��RY餕I�N���}ĖS9���S2L8i�V�"���҄��y$YC��jSM<s,ē�vU�0!����y��,�Ꭺ��\����j�z��Ĥ���e�e��.�ԵkQ���L����;j�� ��@晇��F��e�a;�R����Nz������]��FJ��F>P��qc�W@�!dl9!R��=M�����j��;b�b���a����ژ�4a���jNS�r�t��M��x8?Ou�J�����܌,��*���1��b0�[��?��m`~a��͌dL�a˒�r!?F*
��9x�a)jG!F���	�xt�����JI6��B�OL��;P������t0��ު���H�*��W�$�[��|)w�=e��X��۹h��7���_�%�U���*��PV��'����\��2V�n��t�I���j`�jCQ��4���2�ڟg	�����oB����Ev�Ҽ~#��,�#F�3��l֒��C�Wwxzd'_��Sx���S+�i2� '$N�����ABN:�*Nnݫjܮ�5�����y�=rx����� (i3}�>��E�\Ύl_�j��A0]���|�"�Qyc��zߜ\���g�}��5�X�J�ky��k�E�j�-_Mrc7"5��^�����}�>ĩ����s�<��+Q�R���k�Эߜ�5��A=*�2�#�SS\�!]�g�	��5���"�Mg�W<���ӕ�� ��!�U�&&�.m��X�^D��R^�Z�l(p�cg�x���{��?]E�g���q��-�?�_�Ϛ�AZ�X��[1�����A�F�"$p�;��GBVZ����Y׍���N���h�7�KlK(k2i|x�ħ�A�����()�W�sX}5��٬~�߲s�U ��V9k�s��T�0f%f��(=aU�YYH��v��bwyn>�@s'��pfye��N�.�gFȿu�$���A9��y{^Aʉ� �lzJ������u�Srv@_؝�V'_1n���K��4A,�e,���e�f��_N�E�k�G|��Ow�j"i���X9O���m��!4���w��##���6���0g�#XR��d!w�c�I��/�e���;r�=w�ݵ���/0�C�@&�kP�s���8�x`�u��X�J48X�wCR�莁�Ϸ}�e
�L"R��|���M^8Tw������c��b��������ȝv�X��M�&�j��&i5�u����(zE)���FE�.�IΘ~A�($ѩ��W�Y�s&(�Ҹ�អ�)D���_���YY�*c�ȋ�"}t&���5���H%ߑ���_�����g�<񿰠-�ޜ=�-�\�Q��7�a��EnΚct��;��J�W/�3�����s�<4%VDy�J;a��8"��~v�aA���0ҏ�jjW��(�Ӄ���~A������D�U��\��PG����2�|���.%$#��[j�
zꯄac/^h&ѝ=�Tbf���.�N������Ϧ�)���b_�����h�M�Ql�YΆͤ���d����"�v����^���'�O�C]���K�0|j��QQ5G�������,�6�B/H����G+1�F�#� ,L�0�~���*؏�S|�z���*��	a�C�K��=Y�������0�z m����5���-�Ӏ[�{-�
՜�������_��
mM��A�MqE���P�|*Tp�"z~��h�	��MS春�`�%��P�0�,�\���ڡ�bW��s=��Fv� '(�6?�v���n���D�R� ���.KG�8����WzC��%Ȝ���*�N~�a�U	|���W3Ax���{&�ɋ� �ē���"~����o��N������rz�a"T~3g`|��?�^�$?l�p�k��`���� �!-�%4e-pI/��2�pi(��Cfٱx9R��Q���x��L�-���LT{B�	H�'y|Y#�KY��#��s$0�%�J���噽9�K��d"��-���k���v�)%7`EȮ�
 Wx_�_���v겭tM��Ͼ�%N�":N�t%&����e�cF�(��5b�Z��~r秼e����O�ܐMb�N��ݡt�+�ӎ2����^ O������\08-?��~����IJ�O��2�UKDO��I|���F��{�)I�_֍	�[.��yf�=��GjDnK^^u�<ҹx:��F�v��Ex�y6�j���}�����,]a|Ū҂��-�`k��ǹ�D�EIr�U[ʤ)n�M�I��m�hV����U$qBڴ��ϣuy�s(�@��OE*��	��(4�X^r�x�P�i�?�%��������._�*#�tx���"d_�Z�Pp�g!�$������#����ֺ���0<�C?٨�� c��A���3���i�����uƪ��E���$�8m�ٲZhm��I�q�>=�T�Tm�m�ˢ��;��M���367�
T���3g ��	0�9 �Z�V�gE`�~eF�m�&��2�1#�ﱦ��_�8 )�<��;����[��t�F��'��N��L�d�As�:|/���'���F����p��^��*�uH@xZ�f���i��}�_�`l���ᙞ[/�Ѻ�SBՇkz��������%B�f����S��9��{�
�m�ߠ;?�F�����8$E�q�˘�t��P~!�S�vy�� q��ä_����8x�f\���_�Qtr��{έ`��wI���*�������[[�3ܕ�q�E�>�(�B���N��R�A��%�x�Fo�1Ji7����%l��@פ)k��0�B�g���=4/��T���_x�/�n��,����9zBkG��:ߟҹ�L2Ւ"��r�cb]AV����O׈H����0�>�	��\p`QE���[�UF�T�����nhU��Z�VU2e^)̕��&4(�h�6�h�\��яW�����Ꭼ.!Z|m�cb��T!��ʡ���He���8�f��O5����}d���.�G�|�����	��֩ɹ���A�+��߸]�ں�h�Z,2c���;��թ��-������1��?�H>XBɵ稐�^/�#�9
��_d��� gx&��'���R-$p������Q>K؃�6+dj��f;m�8z_��f?�5�եz�֍KA˄�v;7_��}��nw5�iXs����Ѡ&���	;���X�$:�)C��S�D��j�������S��S׬��� �S�U[�o�
�֡�y��㿒E&�fO����d�<'�-ض�Le4B�}��,�du����׮W*73W
<N&���,Ft|E�۩���G��f�-��8�T�%��P�^�+���$`U��U�1�|}���do�y�~_�3�����ha��nO��>����}���<"�Uv��=��5{B�;���)`C>���^|I5
�̢.m�2s\l��]�@�p���5�Q�$����d0#�PT�*D�h{���t]�I�"$������Ơ��E�W��D!d��F�ct���z��̀�@|��uȖN�>�8^��O�qa��_�4l�m���={T��p� ��#AOt�S΍��2��� �<U�X�k���LH�}��\�
���Hm5���	-�4F���t5��&����SpDUgL�C�c�r`tX�(!�d��;�Q90��w�X�K��PT��=�ĎH���00`�d>`D䚭�$�L'A���w��ES����h�H��8����F��0w}�|j����Jֶ�=uY���4��O4�d�_�`�;��֋9����T:�)!K��-�'+7��>����OWǮ�]�]�袕&&�0���q���"�!NTanF��M�@,���"�3Xx��O�
�UG��r�|�@�Îr�W)e�͞�`�	R��e_&n�I�G�Q���o�\���7���z k48���b_�ui8;���*�������z����qG�踜G�N��'���J���8�l��7�*�{���s���	S�y*�>"H�.��ޘ����/����`���"�)��U!��]?U��G0�Vw+8<s�L�OF��B�tW����!B_f��P ���a��|��J����\��5󦠽�23�0ݺ�I>U�d틽&�86�;H���1��7��^%�黠�7e�����KCσG��YA�����鷜���fο1hZ�_��e��� �(���P����ǽ���x�8it�~��k�fv_(��C�|B�w��'ȗJTHFB�v�E�7*u�s��*;,`_%9�߇�v��x)�O �MkX�=	�, eH�8�JX���0 �	 ;�@�/��4��`�
~%�'z�]�!{�*��u�*q�jeu,�)&@"����y�H���臚��UO��F˽�r�T�i��q�]з�q)�8�,�Hp���"��-󝄚$9�l���-�ߌkBH���M������:~�Sdq2�Nn[���%'E���>�^��ʎ�d�E93~y��|�%Ձ��]��A�����y��� �	���fK'ƪƅ�&�Es�Ek`�L�R=CV:K��bX����8W����Y3"�K��-�F�H%�3@5�%��*�&i�n�Bc�MM'�Yh�}&)��!Bp�������9���dN�ˎl�`���n�!�B�:9p�%RPrD� �v���$3/N�����ƌ�7���AvB'� jT.:.p�ni�ʮ&�J��e1��(�,�
�5V$E4��M2��/D����9t��9�Z�٩8	')�`�u�֯ ���`m
iyW .�z,��jr+@`��?s��.zzܭd���Ц�S&*6��Rp���,Z�㧊���z�[���H�I�,,a(��M!l���y�p�e��t8N�um�<m�Źi5�UdZrM�)�i#���ɘ�������9V�]`�'���O����zg��Ǐhw�(�R�L��h��9w�B�E|}%��}k6�;�=��1=�=U_��p�b��tAeX�����&����X���	��Q��~]-��Q*�6����{GR����Fp�Ct�c����sUb}W�w��721�9'�Y�>�?��$U
e� b�7�|��M���I#�;(�����e(eX9���m��!�M��E���&��	2�/ Om6�u'��Q�<���bB�{%ueC_�gSG1,2��h���[�x ֩l~��BÔrB-gR��:x�F�T������_��mB��?a����S��'��7��lȐBu�y��/�!��g�j���*�YP����B��A���{�:v(E5�#�<J���W�C�Wub���hd���33s���#�Ɩ���{����Ym�]�8a�<�$BM���������g4����`͵��0�rZ�$�#t&����;�y��?iJ��j(�	T�أ��X.�#h�	����F���6�~lW����ܛ{��"0NL�/O� �ڢ���2�o�9ZV1Nn���@\��2	�Ѻ�H6}y<i�_�ݣ���E�f����b*\i�$Z�n���R]���2��!"�H�z�z�[��(�X��BH��#D��<���.�����{0n:Ne�{����Z;}�;�R�0`��/g�c��!����_k�� ���SJ���_u�ٶ�UN��ą��j���|�xk�o��[��u�a��HXR�#M���|I���#�z�Bd�M���;1(=K�bǴJ��	�Uyyt�O{6+��K����ZKD���0��w_\s�:C%a�S��Dt����P1�o� �|�ȷ }�:uynג7,o(�t��A'n��0�:TQpD�M���
u}�xY���ȫ�ba��ۤ�4���~���Ŀc��0	"��N��Ky�f!����u�"?3-���}^ZhM.��!���(��_�W�JÎ�C>�������q�jŗ���b�V�m���-��QP��<��~� t�M�Y[�����}�et(��x�(Fg]�|�UNa���tD��:%?��<��y��5����я���9qu�0+�|�L�ϖ��h�.�׏�����2m�*�{g3
u/��]�c~�w���2��y�;��v�7d�ms ���=/X�u7Ѝ?{]kdPc�f���7	a��x����w93�zr�L^���}�����=���sO�����{�(��xM���F�� n���:F��&af��@:�k� ��5ŋ/�!��什��s!�9)���3Rwe�]�^0�*��Dc���ND���X��J������?D��'5&�T؊� ��_N"g����k�Y)[����Hu�V��,���(��U������c"���^RxA����x�"�N���.��٧���F�����-]����>�+�<2�ӽ+���(H�g��ш] ;��E��������[R��c庶�(��������\;1��U��L�!i��J\���	L�b:?�<	�`����5�i�h!���g�T����Q��}j�d�ݜ�S^��2�(uN�EO��˾b��@^�|I���%�ѻoA_e�%�;���?:�g���]N%�ס-��؜���l�oM�]N��ݟ��4�@�Nk�l��e���#7|&E�+:ʮ8c�{n��n˄l�*ݣ~
�2����I)D�`K�۫�6G�?��X��Mn��� ���<ޱ�&��gċ��k�����VÚ�GF�Q��b�0�x�R�gA6��9��R���X���P
)-koX6U���`�#��� ��J���]�X�@���^�cKW �U}���H��Nre�@+z�_c����K楺������M�+`5����~�5>(4�=�ڍ�@i�/�}?o��cv)_�ۚS�I)(�����|_��E�����ȑ>�8k��\�_�VF��s�(%~���c4(F�ثJ��x|�Z1g��d&C���W�K*��10<h�:�*�4�C��A�G�`��%�c�e>��@� )@��D�	�����ĕn��ê����+œ�Sf�(�fTƖHYx7Ί�3`���RZ%��ap���kJ�N/(��dF�R|+l��#P+�no둛PC-[<j�D���� G=�߲o����/���O���J�p+)^��x�r���݉�Kv��@V�$�ej�,F,gN���xrt�9_¹^�WI�����9؉H�:���W���Bs�,8t`b>���1��L���K�X��j���M�����m2tޙ���p���Tw�ؖ�D��L�W�ד`�D�>��AT{��#C�R��U���W#�jb���$��U^lX��Y��`a����!fb��2�g�$���.�=��jT���p���(((MD�y
bJ-'�_&���^Q���jITd�9B���b�.�0�3\�n�&S��2�EmN٨��o�ՌM���<�}p�Iz�<�p�zf��cRO^:{��viS���ŉ9�/Q��1�^��ry��%��y���NQӎ�r����^�5[c^�"�"n�������]� ![��/�X:m�w�pu���]���	�M�2��́��G���]���g�Qm�pI�+`NAi0't��*#Gv~X����jc&��H��Ԝ���^�s��H���UK^Z��TU��y@���@S W��V^u��pk(a�@��,��d/[`u� �=�����aH@W�7����g��9o��*=��~M�i����%���z<�M��q�r�~�fm��U_)G_T�����.
p]Lt(聆 u<���b���Z�s-c֩R�$j�������@���?��L�}��XPp�G�[��a��U%$2��I�e�Q�*�aA��W*�Y����K��X�9��U�VVU�3���+�é\�&�dW��2�(ӵ��a�-��x}{�#~��U�
�F���\�z?�ُ:y�+"���!�[CwA���z�i��h!f�f��3���W��^�]��R�[)�dT�y��
EC�����HO��.&{�dF>kӲ#�^Pj�"�����X��R�<^m��UC���o�Ǩ��kwA��Q'�N�հXP�^��g�[���3����]�KJБix|�K� ����J�zʽ�{�@��E���e�l���
(�f�qfa0�/iB��ƺgiHme��e�
[	�~��0��
 �N��ysъ����_K�.�������A�]�G���E-4x�QY
 ��Л^�~���*y�žĄl�:�i�1�U^�/�x�xP��%=Z#Ӛ, ��Il��du��~D���5jN�Zś0� ��b�����bu��sZ
w�<ŖIl�WZG1����Y�5rۃ�E0�A�b���NШ�1䏗��U�cdH���-Qvv*C}}`�>k�)�x�.�q>!GǭO��EP:ǉLQ�Y�3�+���5
!�x%���rv���ykr%��5r�K�
��%ů4-`O�� ���O��<MEb���ּY4PǛ�W+�Fr�b����V1�d��d�ŕ)VvsΠ�{����{�o��L5��o淬��#��;:�ycq\A�>=v�ǑXS>1E�T��oW@0�`P�jv���|�Cm���Q:dT,��М�j����^�y� j��y���7���
�:b����ي���Z:�綹 
t���љ��d�п((QKT(17��D�����G�l�Җ��;�-L��.���x��]�g?5QV��}N���eQ�kYt	P���ץ�	Ё���3�"]���z��r^�����oHM �S2З9!<;����N���>#�&JBx�r�^����o�F𓍲`�,�s�����C��.8���m$7�Pii�HSj�W��(a�;qT_{I�ڇ�2W�S(Fa�5lJ��!t~m�O��e�]X�^�%���-��\�&����Z��^xP�b�m�G��!L�1�)z>'/`r�)�]����j5���:b�U2k�b�����`9t�mRy͊A鴩���M�D�#2���.���L�][�g4:U<c�Y=���o,�D���30�V�5z@�Mvs����i{O����גl$�t=q��'`-�ZL��C���̥K�k�j�7W�9���ɽ�����v�&���A����M�73F�Bs�cw(G���p{�/|�D9N��8�[���Z�C晣�W��P��n?�ޜ޽�FA�6���ՉM-��r�|���jn����s�d�������z�7^g$齃Vnի�[�R!��I8��D�S�;>�b�H���2��[��
�F�H�K��b0��4�<(S fb��a�=�����Kiʻٍ�ov�?yq��3r�'?#���OF�gUgT�:ѻ�i�� 9�H�+9��Zm���^�\�����u�
b���
�Yx>��&���̯�縈���~@,w��v�RVnΑ��� I�"�Xqʜ(�;[1Ǘ��ڌ�:a�]��ۇ9g�1�
=Z��t��a�*��|ޫ��S��r�y���q��Z�tF9�voc��K�o������xm�cDD
G�Kε�a�Q�G���%n|w%0fy�O�^�ƈ�pu )g��E��wܽ)�f��$���K�K��rD+������qG�!Y��џ&U�����o�z��O�}A.�{�T�Bi��S=�;�c*��m��'>���R��Rtk�r�-�ȯ��װ���'p�~�x�axY��_�]{�6�Ɲ���ƘT ݀�MBhҠ6�U�q\���? @��x�J+d�cUPf�{p����[��\D�X0
�_=�86�� ��o$���.�n���@�����ET��g/��������Ѷ�,�٪q��%����'N�n�.�W���r�#�i��� K=�Zh�����ʕ�r�m\��
�,�R��1��f���en�:�gC����K��缵]hY1��$W���)N$��D��Ej����t
Ǘ
&��E6q��V�(�.�eߡ+����e��OH�懅6<���fq����ٹ�x�3{�[���.EIp��.������2.�k��t��"�&�х��v�#
&�@���UQ
�^Z�l�'�o�YL��R���Ǖ���� a�9�e撽@��k�@�3��*ɅPV@�.@q��`Z��gc��w;V�eJ��6!��}ȱIy@l&�X����^5���/Ӕ�ySc
`��1#��?�Ÿ^ ������b
@A^�-tU� ՞�)ܖa1��u��`�����P��X�C]=��`_ף���9���Šw�s3�#P�sm�pL�`�aJ�/N��b�(�uMUd��r�P�ԡ��'x�L����	؋@��a��A��|[�U>�AV�y<���{���6����ڄ�D���`�����gu�^�0?Z���I� �d��;obc�S`'��l6�`@�"C1S�l��T:߼9	0]�Y�&jŶ���Th;�r��#qq���]�h��������$ x������,�Z��P���.e4)^���i��t\��Ůt�~}�eA��wRtF��%)9�׷JQ��K�y���J��
�p.�D���t7�Қ���'͝8��kI��ŉs��������ԁ�	]�At�8��Y�@�&dl�U�;껁� (�����*6�zУ��g���û���TA�����h��i1��3z� �4Ĕʈ�`n\��M��6�	/���5�3�&ZCߘ ��v~�t�mwe�6��PI�:�J��P���1���G�s��k�I6�i�2a�?F�.�=:/\�Ėvl)h�Ui\�&y�Z�/����8d�,��ѐ�R�8�����SZ��8��E������T,�GI��ʆ`ĥ�{�&�������$<$ݹ�
�����)��̌.�o�0�V?qy�Z�nC����%s��5��)e�)W�	�X�+b�5����9��"?o�f����,�:L̬�<�s�E0Q�%qb�@�))]��,t �Vb&:"ʾ�{�C6��`G-����m|� ��lh��$$�,�ǒ��tX��jsc�I
f�p����+�i��Px$
M��
<�[t�����9﮴R*OE�T����c-�K�[awP3����V:����?oL�h�)�w��h�<����Z��Q��a�"�H�S�]�l-��=�8�CG�~
q�
*�q�l�dź����fs����}�jl���.}���w��\{�ͣ�hS ��)����f�e�56q���c|�0w�K���I�&���)��/�9 ;υ�h�!�ٯ��`N*V	�wxn�����?FkI�8'*��ݤ����x������5$�Z���n���t�Q�f��`������8`�B*#ݒ[����װ:<�u?+ݛƽ`�I���hD�ʐc�'klu=˞B�mVZ�(7l�iǑ��-�@ם
�wq�ɓc����0+�Sס�9�����.Q��Sz�w'a��bs��6�slw�<g��on����v���V˃Oέ�h����W���
�&��McAJ�oP�a��ƪ4w�;(~8U�7DpG?3��x1pK�_�h������2&Lz���U�=����h՟��e*��?b�����[2=Hc�T}H#x���3MR,�<jzU��Ÿ��a=:�J�D���dR��TΟm1�%'lKP&9�����~�-kP�-ғd�#�-D�+9'��˂O;e���Mùq�3�EU5"��;�1����7܊���Fy�ˆL�Cor�	�^�������a����j�@��W�J}ݢԔ�)��b�;�Ex���;��X'S#�? 0wp.�WBN�c�Q���|��f�w'�p��`v��؆�z�m�>�����*D˕7i��:�݀���ij!x] �����*x���ȳ�wmX 
 �m�<d#���,b�I�۳�n�dr-7�NUY�:�؆�/O�h�������z2g�\R�M�2���)�#�^���F$=t4y� ~UV4���{�mv{�բ[LB���12����(��6�H{��J,���Y�U�z)Q~KNԿy���]Z� �؈�X����R��r��2���Y�Òb��,9z���� ]���Ix��h8��*8#�KF#�0����_��_��$�L�W��.����v9������K���nIB����iw���0�K�v�b�Ř�d�_�q]`�qJ�ڗpp�K�>�#A�Y�1���zu�KT��o`�YT�9��K�^�tT;-�1�S��U.&�q�/���-$�+���d�-F���n�� A�&�ò;Vb��2���xCw*��9�=jV�c�u������s%�����Yk˰V�Zw���*#a;uLΊF���1��[�@�F��c���"�C��zG{���$B��%n����?�x Z�h ���vɔtZ������ܝ>��t�]�D\CG�(��	0��b#٢�{ֱy���5��y �	�Ⱦg�!��.}��͍�<�w���{5ｷ�,�� ]ɻJv�x��S��ϵ=�^r���, �����"o����Jk�?���#j���vB�Ʋ�PkMY�T�n�J@����� ���d �uee���Ж��u{�F=��+s$���Q��6���s��MÈ:�
�.���Y?�!0u��w�f�'���Q�k�u ��."�Y�.Ȩ��}�x�ƍ2*Y��'Y;;��o���u�07B0D�5�	���\�g�{'��~���*z/U���K
�����J�T������<�)�;��H~�������S��4�䱗Irec�FP$9�7	���Q~��IIR�07��b�q��q{JjB8F����w�@�� GZ|-�N"�4-��K��S�4<�Ҍs'��}p��1�/�2o� *2����n����Nb�syح�!ir����";
��h�bsPAe�1�6�� L����ʹ���ў���>��e��O��jj8?b5��~���H���� G��WX�*+}Һ}c߸��l��w�ղ�������C�٭�C	�ͩ�sJ��`]��lEp��)?�>e����D )_u*X��=*H��.���e(�eA��5F�ڭ`Q����~t�W;n��o�U��M�t���ł��92pY�>`*���O��Q
>y���1|�o,ok�qI	A�������82,�M���y��t6���΂�n�`�K����n�Z{��Q�Cm��,���/�N�
Zȧi���Ҏ�+�Ҧ�u��vYFŤ�K~�www.���C避c�Af��E�8P���Ƞ���=.r�A��)$����4ܑiT/z?��u���ؾ ����g)��?.�0z"�NA}?wY���#����
��g����F���sJͲ,���<epq��^��5]�JE�"��c�}� wX��Ũ�U� �q�֕C�#���C�k{aZ,�ҹ��YWE�����IU�Ŵ��E�%L���I\��-}����}FRR�Z1��I/�iE��_��V�"�r�7���A*��c���7��cp�r�:-~���F������Q!	�h��3lJ�..��cW65$-�A>�k�����k�ԏO��c-w%��|������aJI�K]�4;��cq�� ��L�K�	5�a��O\og�ٸ�p?����!�s4��5�y�JU>�df��f�["�AqH���T�=/XO����Ka��K1���h8}���O°�6��=�Xt'��oΝ� �����P)bS�p�.�KT��^���%C�a"zR�h����t�pU�1gS�!�/�G����Um|���!�����}�)��D��E���t�v
�?)S��� ���L)�<N�{�5!,�](v��Lf���3/JV0[��o/ �u������$�8�t2k
uQ�B�ڥ6��l�R%�Ű'��.��6�)�1͕������|����r��ye�z�D_%F����P�_���X�����ϋ�����<���vD����Oɺ�������џ���L�� `_N"[vE��E��kꡈ����}t)[ ���,w7�m�F@�Ȋ-Q��p~���������}�w���P�
Y�Xs[!
�'��{J�Jy�bJ���a=��,X^�V�l= ��QJ�]�?�M����A<γ.�'F	ik$��$�A��"�écc�s��d�
��vHRK>��P�~�X����tw|^�`�e'��TQ�_i����g�A�`U;��ٮ�2�^�AB��^ K�� �3F9U!���h\��9=Ȭ���vJp��\O��V�dBc�v����s�����F�����u���cL����/�8�6�G����`�F7u�,�ア~����v���3T[O`��'ۥ�c�%��-��7x!&	�,���. �<�5��7��D��Nq����S1�ý�����Q�0���
~�ӄb>�M>d��묝Av�[�������ָ��f�Q�T�A�.�<!�"�1Y ,�t��߾_`D@�#�E�mR���Y`x{�֮!�h=kE=����y8x1�g�v�y���(&�۞9��u��u�"o��}�צ��N'�է
��0�����uw��kMҸ)��c��.�4�屏����͓%�LF�V�(Ğ�0V*�l�o'�C$�.*V_��.rU�vӶ�̀�5�y��GL�"uo2���'��o������0���I�n���2&�	^GЫ����V�$E��~ZJ_�A��̋�/�lŰ���|��h�/9��[=ģ��F/4���4����1�CS@���l��! �l���c�M\%V���a�^�J�>T��O����Oԧ�,:�8���C�؅�������T��4-8X!^9
����b�	z�}�JF�1���X�ØM�����GHY;��|Ȝ8A8{��S��\�6��@���U��.�.�*'��{@E��w��]�"Q����*(J1���㝂��_��G��(=����	�D��
�m�<�MHD����،հ�O�ȣ�Rʾ.c)ٹ1ǖX~������Q�-zߩ�SES��z��Tt)%�f��:�&��`*�8>��	L����|��;ލP�V��z� ^ɡ:���ݶ���Һ��@�d_&�`Zg����M���;�4�r��m�|��>� 1����Pa�C+�bW�B��\wS�l��׶9^ qh�	��3�y��v�m��@!�'~��!���4�F�of:?:j�<$Fz)��e��%���ݭ:�����8.
ng�2�Aʦ�SyY�7�'�Y,��D&�FF�j� �����k3)���*�F4y� -E��>�W��8�(.r��ƇL.�~.����h�M 7���P�<�b���7�{S���_���gg�v��<O6�e��3��w\^�l'N9�g;hr����ߍe=�`AṄ������z��a��O�k��ܢ����ҵ:��k�ɝ,��J�h7Qns� �z7��D.4́�Y��*�2a�S�_�S�$����J��3/��i����V���!�2>�5�X�ر�a��,��!����s�MS���c��Z'�T�a�S�w���V�}�R���:�_?1х��?k"����g,����Q]L>>���I��/���N%ͧ��Ąf�uK,	�55�C��]�����8�A����J�bㆰ��k�w�nD1��h&~If�J��}s-
��6(,*2���H1uY�F���(J�;融��A��l��x����f �uS�z)F��8>c��ba�>��%���8��$�(��p8��,��:-gԤ|�WIRi%�x��ɤ^��]�S�o�ע-ćp%��w�O�r� �q��+ۣ�SіI��)�6�����q���
(����%�! Bu�m���0�]=U>7*,y<q�&��a�t�y�����k~"L{{F���gԺ�x�څwak꣖���&rĆ�Ң���oGI$G?���K	���Lh�=��gU��jD��X���(�� �Uo_�����萆7�c,c�'0\�+��H<sA�?�q���r@.�����w���n�>2  �Ԑ��~��B@W�e�k�y0����]px���d�v3�5���p��ߡ|$�������b���,�?�>��b#�������bIi����1�i����S�ܢg*Q�k��~����N5Jc�w�M8�A+b��q�K��`�lp�ڣM��Pq�'�:'�7���9�]�	�%�k����~�턩�2�`x���\7�l�����V�J��=A�{	Q1#dG׷!O�WX@v;^���UXE<(���V(���H���;%��L�_��HO��I,,2����y�k2�������	����0��z�ͷ��G�㊔�!��7h��DV�a�՘�,ʀ�jPZ��t���0x�y#n�V�S;��8��hF��W�͊X�����3@��7=b�X���/:{��9���n;�}U�J�e��g�rjηH��2I��K�TK��.��K�u���b��ȫ�eh�#�)6���I-�8��������ǁ,���W��=�߰1���nDuO���kA!�D���2O55a�_)J!�����Y��¯�l�G敀��ŪLQa7�X$Jܟ@뇜����&�U�!.;;0�g_��kH1��p��Nu�_h���MX�7�b[�����39"�O�d�6�W(�����b�*x� �,�*�m� ����H$���s���*nS.�F��ʨ]=O��;�A1���	�'��j�D�C���7��`���O�Dѣ�o"w=f�e+:�&p�[d<���=�Ⱦ�^��0�N.����A �<iL�t/+Chţ���Ĉ`R���e�G�2����!n1�b$����Do��mZA��z�ł/2R�:H����׏��H���\���t��mm�?�Xy8�	��6��d.����H���CN��4#�BR_8N�e�X�%��Z�ȗ��"Tg�/�6�C$� ]��X0�b�W��l�Ȓ/�Jj����������oI^��h�b��{ɼ�5��y�q��,#}9>h��=g­J�M�ʉZ�'��xA\$&��>��mM0��@��EAjzR,6 �H9�	���#՚r�`ݥ}3�莠������� �� �~��Vn�1���:6�}~E�Km���īpC�m �E'���������wjd9������јW]���,��2jk���9����XL������kkrԶ�/�U�g����K�$�٦�/�J�䩦w�y8��ac>I�==-4t�hm�ҕ�Tz �<�|�f�e�MN8�I�,/9�����6��e*��`Ѡ*J���e�CU�Q���Q)B�����,����h�j-� ��.��ۿI�ADRC�Aڴ�X��6�mۅ��$�%��*4�~
<g�U�f��E�}=D5D��>E�����9��C3"�r��.A�3�:����v����L�zŀ�>�I��T�D��>�R��$�ym��0jc����E=z�M.=Kq�0�JT�D*�Ù:6��W-���˄�Z��O�Sm[�4���
�!8��i+�_�-ʘ�ml�Qf����[r�ʚ4��!Heg�_lX�B�?~��7�+K�r�
7i��54�}C/g��>�{(ۇ� _�8֛�9/�9�ڲb`_&��O�d=H-��U�z�2�r��#��ûD[������cO/
V"�B'���=9#ˬ�{f�-�u�rH�s$D���K��%�L�,��6|! Rk{�`�L��3j�;$g��AAWT�Ͷ-E�2�wx>��(��u�g6�3���}(��u��`�Օ��s�g]WN�K?�q 9����x�iC>;�vy+,��`(�CR�5
���w>�Y8�3��6H�;��lVZ`�3�`�xOV� �8�k$_�\�`��1Y�����pgY�>����w��&\^~-�Q���eA�׋x���(��H�	9��7Ks����!�#dvv���
D���62_�"��ꎲK]�v��zH��e
��j�= <S1�~�MOJ�B�C��D�v(�H�S1�  _���\�W�^oJ�<�>1/��GMv�Z��cͭ�|Xr�;@V�\���&�V�Je����5Ԡ��=�1�jX�Ȧ�@�KP8�*7@͊~����������$�"h�T�~α����Y�S��Ƕ���ܠ�q�kaE���2q������!P�8����\��8퓦Z>�y
R�b�ʪ.Bc(~ �����$�J{�[,����0˪Fǧ6�<f�'SN������NU&L�7>+��wi�ةS��&C3P&��[�`��錹,a]kBӑҾ�P�p�}5g��Jz�U9�&$=�4P{X���1J��Br\>�ɣǳ�����m�e���ۚҦ _�.�:�sk�6��e=��~L�la�Q^�����Y1�N%�n|�I���`%ǋ's�*AL���A���ON��Va�����%#6��el�d,���)	�ʣ4`<-��L`�sa}h�C�?����k����;O�5��=+{�
���X�7%��71�MʓconSl���(����l�u��|^E�֗wm� X����0�(�0����-8�-+w�ӥ��29�AII�A����"1�lA9B��k�>'���� ��;-2�}Z�fՇyǌ�{H�6O��d�P[]l5Ml�h�z��.��yw~	u�sGt�������p�m"����	������T�cD(�6%*g)$l�n�
�H���Y鳼D�UѯH��%y���9_LZ�>u�^BGoM%K^鳎��@��G�+,nN��B�v�X���`fGD$�=<�Y�I��K.�Iu�U>��*��օSC�Z������,(}D7�1Z+�W����+��c�qZJ#���-��-� ���OU_M�����̯�ַ�C	�\�>��Ћ�j^/�^rel�h)0zʳT<�zi��d��;��J�%��� |!j|�4�] kpEʥ��Cf�IB_r�9=o5��Hh�3x;��F.����$-b� Q���!�'<�Tje��ɜ��妒]���qAWI�1��B�)ۈ��z�єd�-ڌ��+)(�E��r0�9��@X,�o���-3'���UӤf�{�*V�u؇��'3oߏ�2@�)n֟�>=W g�}�X�ԑ�|��/ϴTB��z�3��])���-�cd�R�e9&�LDb˳���!3������7�Ea�f�F��s(3�G�xY��?����$YHF����+e��~a��%���2�8%��6*����;�J������4Ð*�)�!��@���ÔW�y쒗�>D/�u�2�9���\��f�v$X4@�ĉ��:�S�m,)���
�=[��NW����;�/���Z��ٞ3�������d���2�0�
�.����[&j��GyE�G�U�UK����~�c�w��P�,sK�^A���>HpT,|��W֖���06�A�a��`�!y�>T#c��QN&U�$o;c���a�[�
<��*) t]m�OzO-��������	�[ZDm�!�E�^*ҵ2	��_��O���e����Y��V6��m�7�s��`���o���� �Cn����c>�ꂚ����0�9�	���s��2�56�2Vі=F���&��]	Re�4p�U��$"�=��j�čO�����t�(O}���o����m�~�,�a�l]a�l��Q[�*1������,����=�1�̍����z5�����F�<�~�D����3����.�n�fҐz�{q� &��`��W��Z�o<�/�3�HC��76���=+%i4eJ�$��~P9�1	Z�װ�9[�,x�o���)�%ش��p������UV�5M\#��s$|���e;����1o���*E
qh9�Ys��F�4����Œ=]I�e���@T�C�F"h�����qS֒G����*��Vd�r�R�����7y�V@7��(nB��u���W��F�B��Sh�&V�*����d���7�o ��X�L?-R��a\xr<ܫ�]�hEjl4
]>.
bh����7PI��Ua6p��wb��r�=&/������>����2Ѳ5���>t#F�a:�[�s���0v�]k^W�����p&G�[� )�q�r�|��+ܘ��O�5Bsh�>�ǌ������<��=n�[t�{/��Dp�ƶ�E3E��
��~�O�щ}����H���";}x���/8��P�|uzC�C��a�bI����N0LS=���#c]ԩ�f��Y.i�k���ફ��(V�8o����Ztc�؇�y	�ɲt�>�-�vi������DS����`�YjNxrZr��t�k�r'*F��K]G/�+�ݓM�>�yI}��M�_3�*���[U(������zηސ��h>e;ٙ��_�V/���5����r�x��&묵�
���B&Z߈�z��[�z�3��-V�. :������-s�Y�t��Kv^:# r��Bo_�{M^Ģ���2	��b��BS�-�M�M�
���FT*���eȲ4�j�s{	��y��w����Q.�tX)E�'ҭ�2��M�/Z�.t��<��P���X	D�矾�)n��[BK���� #Ι6n�Cz�L�~9o�0]�=?��ų�,+&��g���buSm��,��r��ko �`4�u�%O���%Rkf1���V�>��8������:)�VwCq����a��2��U��n� ��`��7:�\�KG��Hi:���Xphw:���9n�R᤺�.$���t�>�������Ha_ۢg>�}����I�3�aI������Ѡ�bv���:�N� ��:�y��T@�ۧ��F���"H��L�I���D�9"����s[�&�}����$�_�}m���T����Y�+�V�nYAk�1�kw/=��$J\��+h���؊��WBo���2[��b��Te�*��$$Ѹ����^V����B"�=|�/=q��i���������$�1j#7�%�_D���蘒�%v�o��XF8u� U�s���"g�[�i{Ǯ2M�s�uV��Tf݆O�����m�}��W���!���Qt���d|ċ<#8�#�_�d ꃗEꂘ7<�	�㟭�q�c��F��y˥��/	�Җ�HEsE��4�[]��h�d�N���D��)��#WS�ƥ�8�O�y��13����[�e�wy?���i�gA��9F@버�X'�9��\�����=�6�{1�D��ScT���KNԎqtkӐ�%.I��Z"3#���${�c��ѿq���õ�g'�(��9���cˌH��7�Fg�4��ANS����o ~�IĞ�?F���6�)X���v��EN���*n��˥���N����5�(��.L��.������������(t�\�r2\)y������ĳέ<� �ۗ����>�ё�u���L��-vR�q������o:G7:U����TL6��f׽�+e{��SuU�����$|9��A܉Y��9�4!��M*?1x>Q�S\��m?�"�RKIIC�]��ٴFnX}-�JC��f�Gi��+<\o�KBmy �WV�KM[��[?���6��O6���$����rt.�մQZ��l![������:��iUq��@�n�Qm��ne���Ї�i�7���+<�t��IY|����W;*��FG�0;i�xX&�^�O���>'��N�e��s��$n�MZ~�z�h�h�`;RKx4p��{�'�E�6FQ��r�m^p���!<�Xg��I�vs>�=[�����3\|L�so�"����9�E�t+m�Qe*f�#t�ۏ�O��'	��ٕJ����}��Gk�އO��d0{�G6S��܎Mq'Njr���><�O�yP1^ޥ��H�tI]qlb�Hm|���a;�q�c�4���� ��Æ�D�X�S$�Kg�,��������n�ӥ��K.'O~��&���=�#��@�o|�s[д��ΖLl����W�Yo��J�y�F��&/�[��ڣ!-����
Y�G�ioRI���g�_���22|�®�]x�4�:�6�.o�?7"�0@��M|T/� �H/@�X�w�z?��ǵvE{�	�t9$�$z���:u�k�0�|b征�=�;�� &��g�!鯦�'�[�d��VM���;���nH\�L��j�⏯���p����,O��.�:��#��#2%3��u/��u^���[`v���<���w��`|e��*��o��&�6�	ԖW��%zeA�K��y<����R��Ng��wHCf9n���+��H�0���+V_����_�=v ���ź����+O�R{5U��(s�`���9ۨ�k���������H@(1��M�������i��ZԉLj��v\���XvB-I�N	Hd1�*�Zb���x�6���*0]���&֘�b�:�K8�AՈ�p���sg i�6?<r��?�,҉Vߓ᭷pQB)�hM+F�G
dS�Yek+;�e��0�#��}��萋ci�S�\v�42��CP���w�z���2l�r��k<��=��Qq�rns'���������t?����F⑿Ѣ̇�ު����<�/�s� ��	`Ұ�̒>��� ��^A>0hì�ڱvh;6�"�w�Mh��f���	���A�k�q�+R�@z�?Z�T�u��y�G�ӱ�^ ;X�RA	�nѴ�۽�T0��>�W	����Rه��7ET0�";����M��$h�4�}wx���-vRz��>g쭐�[ C6��^Ҍ"[�˪~=���u��������qV�#�e�����k��0�s�hݹ��b�O��7��)�OT�����x��#%�o��.(�|�'�"���T�Z`Ƈ�~���!,.��u���ż%��P�(��۱\Q �ӧ��gδO�=�7Ä����M<�t/a��9F.>�e7�y���wSu���G���k�0u@�;����A{ʉgZ�AE:#��ˀ�~��f�jP- Q�-���>b�/�B"�v�?����r��Jj�:��O_>��W��Tb�lC'�8P�Z��TC"��r����� V �(�z�K傲|�*�����O�z$y)>�P@�2'��pBLL����!:��5	���R�ի��ª*�R�պ
'_~c@�d��l� �f�u�C0<b�t��\�H�x�}^%�S65f��J���R���/q�sAM��>�˱�$P�Ä�[F+۞e�����,��H>�b��֜���~?��-!KwܨC���U5����$m�x	[��t�?�#�<gdC�w,޼�ձ3�������"-&��e\�I�m����:��(_�i�3�:l@E	�����Z �u0��35ZӨ�"�+������S��y�ׅ���g�Ρ�:@�q����O��Ղ0+"O�Y+�h���=�DXԃF0?iq�
�1���U�l+�����Cve�S�Yక���������AгuW�.#�\U��.4h��6��\ p��o�梠#)�����M� l�;�1�E�j� �����UyG$jK���У@j�~���-�,-����~�&m���<�Z�B���cC�rS]͕^���e��@ڲ�=���� s�j"�L���L:ɱ�7<�c^�����r��Qx�՛��ZÇ4��7���	�&���޽^�M�께e*�ɨ�����..�׶�&m��U�B7gY���}�"}9�o��B⸥��~x�w�b�=�b���� #>�9��L���{U�9u�4��6�(`3��הq��6,��y$d��#@�i�D�p���'����W�7k���B����4��ph�?M�M��G���b�hp��tY1������u�}��[��.�l����:N{��!說�� �c��td�&y�X=?G �v �i�2�Ӣ�[����F-�e\�P�"�{	���MX����ކ[���9��RYϞ!���܊̾�*���:���H���<�p�k�2W���l���Xʖ�5�[%O*���n�SQY�Ϭ�E��������bu���,�����'�P0GQ�ߝ2��;�
6ӏ5EJ[U��82o��w)�1����:�qI\x��r��E�<�U*�B@E��=���Zr ��,#�O�U���2�o�`%��p�I��m9OGS,�N�M��,yw(0xO��~f���(�|D�$"�X�!k�UG���"���b� �~�_�F�΃k�2��	�\��#�O�\'��آO�t(�$�j	^P�<��X)��'�-IB�D_��+t)�9�Lk���QQ��XyM����S��9�
؁7`b��;n�J��4g�no��W��γ&\[�=h����E�6�.i�\I����k�l�qەq>a�Dc)�I�P�֜�~NB�����A,���XJ/֔��"\[�]��Q�u�G����5}��G8z����a.a@��������&x=a��5F#�	��nqOGC����#�]��.�^�S���[�\cBb,B���9�#�~յ�ޯ���k\���N�����W����f�B�Hk����QN��8��_���Nד�0{nc��#l)zo`<�h��J�ձ�>U*����r�Ҵ���m,�9j� ��E�Y��%�,���QQ��ǟ ��2�/K�Հ��T��0�A��,����}�s�i�佹����tڪ ��v��<�2�bp�a&�p���Z͎}�`?��'l��gh�G?,?�(�i�+T	��7��3]��'�;b�#��8�v������lU�Mq�\�X����ވ��8<21���$sE��_oy9�u���f!N(�kO�%�y2���2qUPyd#1r�A�R_pN��Y�Ҏ����� K�vW3w���ե/� E�2�G�`�}��4ߙ~����;�v��t�3иgX?A�/6��O��-$Z��T;���I	���d1'�tFSsv�z S�d���ja(��R<��[ ��6ջz��d����jX��~۰Bw��>����i⩜x���bI���^ܖL�7�i_=gN�� ӳf�{�;N������k��Q�i�b��);0�C����m���I��@EF[6�{�5T]�Z�Ёw��;UR�)�"O�kc��1?��EB���:�dZ�1����� �e^]i���}e�?�D�˥PP.�s�na�~tOW���]B��۲��ߥ̱ufr�c��٥���7,�����ixc��l�H��W�붐�륎�C%\�b��G�m)���W	�s��}�0�n�6LI�B��A	^Io&��g�@����;�8?�Ѯi��t��&�)>AD�V�K����Gו/�����тO1\1hz6�/s�6Ѫ�c)�nR[�dv�Q������[�b5����a�uk�k����8�q_5��;��LNh���A� �����'u �W뿀~�ӎ�&�)AL$��l�r��Tړ�y��t����&N�U�[�ͮB�a��G��A��
�ݼ�0E;�, �vک�qH�{e�M�6GZ�����s.�̟�:v�8}:�b-*���H��<�)�+�P�`�a�C��7�'���5������؄3�?p_��V��eP�X�s��]Mc�5���A�k�Fq��U�j�5�o��:B��,��<L��F]��QL���cOk�LuU�e!1�a�@ s�h��^F\� �bޣ���U�\-�����5�̞��˧&�I���O)�B��EuP{M�4�:��#?V�v���צ�k��?)��-92���v���)˴Dlߗx��+���|��3������*91FN����Ȱ�Ʈ��.��
���s�Nok�PQ����+��c�>9^�(	u��Zg�dz���t��Ϡi�q�E���{>S�U�֧��~Hմ�PֽU*8��
R2Y�vMIza1�CIE�-�G��?HB���$:�<��їХ��P2�痌^P�߃��ؾɡ�zC�
� �w�@���VC�<82�G��������r�&���|} ��ٰc�ۿҝ��E�ͭun`��4�+�F�eӨ�YԸ9'g�I����8D�dU"@W�	V�nZ�i_�c���^�D�_��tbC��t��{S��l�'�td�A�\P
!��AP���#�v��"L�\q�t*��91�C��4����"�+��8	��4G� =+�^��&?��VӸʕm:W��Q-�ky;�bu-���
ߦ���R��B�ޞyrM&k���u�)ѩ��ܰ�{x֚�0 ��=�x<��}�a�q��(�~,��'3�yD��H,~�lp�{b���oaO�l>���ޱƫ�?ܶUΕ>؀a��m�,�Sn[���z���`�r�K}���%~.��"�<X���;�o[]������Ut`�Q"�{�o�-���C��ڧ�R�o���5�� Ɓ�LZb�y������D��Q���~���7|`
K�a�1�/��v)-<ک���:�<��o�&�\��h��,��ET��/g8��Lx&���b-O�:�c���
("k<�C�)̕w�w�:�ְ.<_epxZ��R���2�3����Yң*�	J�W�)��vj9�Z����]/�w��O������'n����
�XX-b���z��TP�i��0g�X>Y�[��G�8�V�{:s�\����G�$�e�@�v�L�Ҕ5R������Pw��-�Om��B65�F
\=�:���T�P����` �o�W�%J�����65�уZ��2�_���:Qo��U�P��l�X�ɂ��bI��˹���Z����GA��� ��X��òt�ʅF�j��?��L��q�����;�OF��,����G�g�U"D�{#-�
���;��t�#�[ƯUɓ�O�蹝��C�mD`�粐^^
�f��a䗓��ֱ��$j?cGo�i%�Ǯe���`�n��U����sŭ,
�ۊ.�*��C�!�;$�D�YL���
�u.X��?�\#p��a����cA��z�2eCY��	��?�u�M>p�� S:�$9�D�u�p�V�oɷ!�c��&�ٯ���sԓ�qe*��4R�&�ȧh�b"4��$�J|01�D�6=ez0���J���$�E��1���9o�5�T��o:Ӳ�±��YǬ��o��C�<�p?H��E��˃K��ajG�K#J�#{@�$���*�������G�?#C��3ư�X�݋��?�;5am9GŸ��q�K�Γ�Y�F{,�r�uӒ�yO�Oj����
y�!λ-���&�2�R����\��qo��=���1�q��4�	��QY�m���]4C���f.��W�@�G�&�ZI9N�\6�������~�ϫ������7�Jk����i������h���&�R�`i��.ʅk���E�A	���'씵��L<�9P��N��W�Kg��8{NM ��7e��ë�s��
tb���@f+��;^B^:�F5����	�Y/�D�6қ��8 ����3�л?
]����#0�")�Ǟ��Y)p�v?�_�F�"e�yv-�6�3&ė!�?-�O314v�"C�vҧk��g�"�;p��D���ȳSq��鳩�^����� �T�)g�
�U�;׋\wNމp�R:�J�7��{)�bR�lR۞�֝��a2<dv4zT�匓�Ɔ����	T��@���BZAdpm�p�OL%���A����k���*@Ҡ��ң�q��
B&�μ	��\Fj=�ɞ�םm��| �
�:J׫�C�u�h6���6�WJAKH෯Q0T��͑�x�ET���JBҿ���+���5e�	�{�ۢSn#wæ�E�m0�s�~m��C���:9{�bT}&ۍer�8Nb,��z�O|
�K>T�_�3�c�#��s����	�� v�Ea�bZ��5ˇs���]�X�=-��(�!<3�t���t|�5�&���^D����	�v�Y;#$�/�wI��9������l���ƚך(��ׅ���Ƃnś���>�띨��������>�͋�[# ���l�����*�)��� ���7�-��(�FS������l�7V�}�4 "bT~�+B_;��M�f�(�j \�B6"cD!��3���{�0v�P`��"��0Fn#R�9��y�(�
�:�0q�M|j���kY�B���)�)��d�pg-��؞�ei�&E�T%}Ys-��H�RA0�mV�kHC��^�:Ik�;H�Yl�ƞ��Tޙ�O�( ���J�!��-���x��Q�r	X廑� �j����a;��8������$9���裟zDMi�p�W�w�����i�瀯�V��+��E�ۚ�3��q��τ`l[�~ p'�}�"�� �T�� 11�9���w��G����u���l��洰�6x��Y{��Tk�r�j5G�pwq�.��-3R��\�ȹ��h2��+ː�Z��"Z���ϻ(���Z��})I���#=�-����]�275Y���T�y�Mf�N����U��cM�~D<���}��A��&W	^�y$˻r�.کӮ����t=��6�2��#u���C�X&ۦ�jI2Ů���p6��"�"��p�ҥ��vWq������
����gC_��rY4���?8Y���B�Ґ#�N�J�L���9˵W	l� Ͳ�F����f���}^��ɇn�J4��o������TxB��'"_'͇eͦ�%~K�O�u��sN���+.o^���A�=�=O������U��0��2]���v����<R��c|��8
�2�b$R��BS%AMJH%��j*0����қ	��s�ƎF�3�'Z���-D���.1���/���>�P��E���!D�Ȥf2�����[[{ D�9�`�L�C0Ҕ���m�G��L�R䀁�ם�E"N;�y��<�F@ZPC�:��U��-���Q�~_`񙟆^�Bxin���`�u
�C���T�����tDXk�yc�|_d�&mb��rwZ�'�:�d�Q�VE~��d�R� bv+ �������er(h^z�� �B:V2Ђ�K�7?�v?^d�g�����'�$�y>;|�1(�ަ��5A���1(�o!b~p.�u.eW��؆�	D�i!�����8�+Ք2I׆�w�U�^�>�<�9*=��/����ݕ6�oES+���e���p�����U�1ꯊ�W0�������O=W�z�c����Z�{H�iɢFF!��F�ʓ2o$���eWL6�Q� ��-as;3|`���;���Q��_;& ��"����d�;!9��s?�`�R��k��M A�!J��M�eF�c�u�pU�MH�����M2"G�,iά��w�>���j8a
 ��S�?��C��LI�b��.�iOm�t�^
ym�_4�Ք����.l`��j�o��$�M�5���K�%Y�6�NЃB�͏\`;B=����@�E�9�yfm&YN?F�<�\#�vY���N��)�Ƚn3o�;�m�*X���AC��Y�s�4o��cv�1�� ��qAzj�n��?W�ʳ?j!��� �!��1{ћa�g�l�AU�h}���Բ�x��hHro�"�W&j�d�5��uedMY~0���xP�u�p��x�B;?�tBL6K�%J�� �өI*�;��M�S��% *�����@�E���������eb_��|[���>�Cf8C�R�ֵZc[�4*�� ��)�'�wjP�\����֩�d�m�%�����:����9�ޏ��4���U�^I�,�UmMc������!x�5�<ڣ3"������u��٫��2�=wr���S�2�@�Y(�� �F�[�9�D���r ���Qབྷ�H~fwetJ�-�O����W��1�v2H���� �cn�����9-n)�+�î�R~Q�����kf���:$0Q#�=��I-����j}$�-L��f���R%��``�L�7gj��?����s|f����}on0Y�)���S�!}蓊)�u�DI:��lO��U�,�4���[��&���<����؂���P����.	��u|H�x� +O$�6b���D���N���0KT`�m��]�M���r��bop=�-��O?�����#�����^p�c�X3��AQ|n�_��oæt�S*�s�C峲4�,���6�/p��P,V q@5��jy��Jλ57��_�9�O��_jZ4�=s=��$K��'^E2���)���E���.���^}�}
����պ�wh�� |�����g��B�$�o-.TP �b���7��)ʞ�+_?��'�u�o�unI϶d�~�m�[Τ6.x�t�,���Q7ab\���H����Y��I����*��|��Q�)�H ��}5rV�"�7;��<$�@��!*J�j3����/u!��ϪiU+��� �JF"O�"</�\e��#�笣,O��K�M�Izf.�.�V��e���)>��͍Ҥ7�> _-���Ġ#��(�)�W	r�]�_1��}B�eOrF�I$��t� �F�%ǻ��Mf��N8���GxÓ�9�ghm���R�
 @="����b�1y��s��+���i��5�#p(W�\�t�nIF:�����kw����������?!�޹#
j�%	l=���,5���5l7V�2� ����E=B���@ �r�����oC�
$�*�Μ�W��O��f*g)n��?�$>�����X�j��D��;��p���a�"�J����i���,W������L�e�/���ks�m=�?�����m�:�ߞ�[��vS�v��PM�f�D<�*�wI2D��'���5�Xˣ��\��S��@�YM���Rه{�q�0W�鿑ls+=�p����-�*�ȫ�:�a�w}�O��t�<zj������g��O3�n�Z�_N��V�￈�H��?�=�wQ*�b.ۨ��O�[Zݦa��.�ff���H�%�f���L(��0?am�|�̈�x���; ��k+��^(K��l�����BN����?��d�w��\)Ƿ�S��s��Nb,��=_w�> ��.l�<����H�h��2�ώ����`vB�&�ߥ��oZQ�K_��xO4|��h16���X�����,ru�a���G�Kbe�W����<8,q
{�Ϧ�s��Xc��n����hxy�ד !ɳj��1%{'�͙�g����^`�&{ ��{$���H4r�@�é�~Pzn����ʭ<Z�@��g��ܲ�L|\9$�fP��?h��wb̊���%v��B��TX�bχ�&ǪrÎ��
ކ"5���@#r��/+nxi�{h:���ͮ�V ����ΨkByu�M+~*�.��}4�K����=.��QԶ���m�K��Sr��?L���8z_�ȶ���*�w[�o��Nt��q���9�I��F�ȟ��}��`ÖD��r���*˸��4R���y�� ��*L��d�u�4h`��?%k����� F'~W�5US��B��~s�F}�:7G�W_
f���׊����up5<u��t���~����#q,+#����o��1%r���n6�t����5q H�|�3J+���0hct�8 Ь�2Y3wB�<=�)[^�w=-X��qY.���!Ç��.� Z�A�R9C(#�=�4g�"򚆻���]���A�t��
�M�b\:I��Ӫ1�b�qJ��`q�RZ~m�^&��AU��9�'w���o"��tR��s���a�zeQ��o�L��<�W�fr��Al���긨�2`��2;Zs�JHq��s��F��r�$�'�w�̤x(}�E���9�� C}w�l� �Ǖп8E��;�D����oόQ�ѥ�D6<6�`xq�a�r+�i�_}��]�� �dOG ؁�P�9_�9���+{n�"Ll2Յ$���Ҽj����@��?~c�e�C��x�L�n�%�E�JxI?b�2rhe�n��X-!�~�ͿKmJc�@��6-G&@�k�RY� %��+���5�G�m���҆�~i}���|�lpwl�1�"����9�PUE����I�E��_,)�g}�hA�K)ҡ���3r��nz0���L��gF$��`F��O�IV� ����5X%t�y�7S�2^��7�)���sUt�^���Q=ݶkd�w�;bB}����|�\�Þ�#�a���$�:�+�IG_�*�Դ�_]d�7Ps�P�n�o���3HߙJLl�h�ծ�w.�_h�D��1�x��$���\hqO��U�M�WM1���q��"�_�OLW�����9S����G������HJފb������g>F���<U��Q�:D�v*�R!�g�<*�<X�٥��{��1-�㷾��ۂF,m�a�F�<Գ�!PG��ޞDhB��E_�?�9��5�c�K�XU\d-�Ja^[yX��s5��JST��'��3J�3�3�Z-]�: �K؊u{��&c�P:bapj|ƴ�Rl����O��y�S�w�鱊����o����@,�g�R����R�5\1���\�����ɂك�UPڻ-���;�g��E��ު�y�9p"���_6�\j�J����>B�`���Q�(��$�	�s40����)�<l��Rg������L}�`������8�q� �}�Z���8��C��{W��6��i���k��SÁf̞C��Q�����ppۑ�%A� 
'��`�>�Y���;�Lz��#H���qPc��ZA.���,*��g�K��ߟ������/<�E��?�j����I��LQ���T�ty1��b!z �\��a|��ۃl�/z�s�Hm����6�t���͞�����QK?�e�)Y�?M�f�t���^]�$��*���gUm2(F��.��ܛ�؄\��.�B�4P�r�^�TL�v�Iz�Ĩ�vC�'g6���>4�oH�?�p4�|����K���׳�h��l�rI���:�z����[�PHX���գ\M#$�<2�9/��rA<�F^�1vҍX?�v:���� Gj!j;��e�z����r������wƹ�Bf����jlH~�]�:�8'`|� oB� ���[+U?Ý���1?TLz��5NUdX��~@K�b��0!$���/�c�e�45X>��W��[˄U��
\:2�ˌ��:z�HR�1R��i���������<����Bٓ~Rd���a�?���@��z�:�z�=a%���c��D|��L��_"}��x�Kt��7���bn5�n��������}�-���Em��{���$�6��V���,�"��8IM�E��6��6�y���;xz2B2<_åL�Y��~��B���RƑ9�p���kĞ�Ed.��m�)):ә/F���Ab_�P��52Z��<ࣨ�JV��J2��5̱����H�d��B��c#U�'��p�Ԝ}@[�[
��%�|��[�[^M�)�c����.��� \�!�D(t� %{cD
��=��S��y��`A�2������W�c���^������G�K��C.�/K���L�_D#�U���q�7c�K38K��1�>�Q��5���!Y
��g�Z�$�y���p�l�.ܙ6��J��/�*箌!��w��(s^�71>9�U|��?�M7� @Q]���W����sJF�� Dl3uo�Q����b�]ޒפ�v^���ˑؙkI�B����
�O1Q�'LK���w�$.ְ�𱾵�$,���mO˗�B�˼������ώ2�,�eR�4�_�˨W�K�M�%G�-�x�_�4��p���M�(y��a9�~�ߋl=f�зmr۟�p�8G��P�������-��N��S�8��Gk䥚gV��xR��H����$d�	r *��`6����]~ �=j���~`�-7���O6 ��B��G��n5�ò�E�ܕ�t4 _��C)R%vI1m�4�Y�������~�fL�zXc߶P�yR�{	Y�L+7�[^�"��9`g%����	����cf���$ô�ᚦY�_?�E�	�F�U̠��~�ʚ�f�[h\ݶk��(>�j�n�<�kr�_|Ȼ�m�+Hh�h��F|��u;��]��\[�&�;:����y�*�~Y��a�(k�@��wJ}6�����*AT�������M���&Q2��[�ICC��߂BD����E���B���ʓ]u5]&#&E�@�U�`4\���Ģ��: ��ꔘ�\ތ��!��Ȃ' �홐��ȓq
;�8�f2�'�$���UQ*i����D���]�N)D��%Eo�eV���q_�\Z��h)5).fqP��kz�a7��<q+��@'WG�ή?��w�U"�"<c�|oZ]�(!�kH��cc��������+A@��'�	�.����X���b��,�<�^��!6;�(3�@.k-�-|v�E��)?V"��i�^�^4���;۴���ag�M˄�pMz���Zf����]����,�P�?J��(�g��:4X�'���Me�� �<)P�����Ag�/=uh���P�f��5\����s�] �rV�;��؆N^�,Ls]ItF�ٕ��"��xL�B�v��a���lۦ�k�k����L��vlĘnǡ*R���$�6d՗u푶<�T�b	\��n'd[pA&w뢜&�I����T�w��/�9\lq|�PʀA�mn�Z}"�\�g��\�՗M)؟L(�)���B�$������kP^V���t�`�2��0��c�����_�h��t��tq��է}�*�Ps�E�K�ϫ����A@��8~F���Q���'�.�E>-���j_8�Z_u�y.;���Kј�&^7�y���ɯ/w]�u4Ο�T�ficmh��h�v֖��Nk,ALcW ��'Y��W:
���l�Fz�9Yn��x�sfG�>��vR�(FG��C��JCpSmnu�᜙�|�\��*:�۞�@�Ze�|�<gX�LNsD0���.�$}&H�U���8)$U)��p\���,�����ID����l��o���H�ɺ���BaԼc��+jQ�Y��C�q�i�sƼV��l��%vPC��I�Zd{��0�Δ�QY �=(���T*�iQd
F:�ݹPe���E�&m�݇�jy�ִ93[����:���)k�ǟ���+�G�P�:�sEL�s��B�w|ũGTgq�!��5�W�eI�ؚ;���oH�̀s^ۜw_%O�eؖ� �]G}��6�o���~��x��|�ˏ4�0����ֲxֶ�Lq�fiW�rA$( M<��?��`�&ȹ8�Ww�J�W�C��$jNy"��q�Ԥ�Q΢�E�9�-�FO""Y�9�&!y&���!,~*��4����� ��~j��~��f�y��ygY��+�4��9���/�Z���r?U ����=>���Z�ޢ��3Ij#��C�� 	W�\��U�\��O�"���Yd�Ё��0[�s%��<�N3A����}�H��VD�F�uQQ�A.�{���+JJa�2l�]�Z���"{���S�
��.V5�����M��g�'-8���V�,���U/9�	��߹��Pz��R��ȴ?�ݰ=�tk�;�IlVeO��t頳���x�W�=D�\rl���L���g��~�`�G��{n��*�S���Γʂ�hI��R�ߢ�����@ݮ��q��|c�������W����ڙ��k��؛rs �s9�(oXTj�mȡ�65�L�Mh�X*=�Sz�n1��DP0��f���Eݭ���O �ݬVcOZ�ѱ�һ����iS��&m�O���<��%n�����J!��EP�_��:+����Ι�a����3�8Ћ�>0���?�O*�mw�FYgS:����{ߑl���'ޟ0��M�p�Aޙ}���I��X�B�m:�Q!���z�R:��5oM�1���e㺧�?,��S������4` ��ږȜ��\�� ED�ܸ�W\������a4n��ΖQ���#�%LӲ��aK}�*���@Jd��Xy���1v���Tl7��421���+�&LI�6Ɓ��ت���A��T:�"V�*W�˲�:�[yE�n�a�x��b
2���9P����P@V�.���^P��G��9�M����Z����5�+@d���ju���A6Oڃ�hƲHܴ|J���`lj5��T��ť!-�h"� �د�Vƭ���&�� *3�H"=h}ƃz!��	}=�U�8J�/W�D=n�ؙ��֒�d
n�<ړ�"�.Z9\���'��Y	��j�1���{��N���N� |��)���������\$�>�HV��S��D�aP��K{�3&]uk� �~ET\F�'��F+�m�b�*ٻJ�C�GY����0F *R���[[�'XMp\�w3�G�荦cS��b1=�+۴��z�?��1���*��/
1=R�I#�2ֹ�1l���$�]'*72)�3���..O���0%�at6�ƁS�N�;o��v�7�ߘ�@�������Ԙ���]���EK"��b��%[>����n/ 뚨3$RÏ�m}	qz�1E��'䏒{���P�#1I6�>��W:?�F�\�!ݩ~$��R�o'e����K���"v�<���a���r�'H��y���v(Me�@�S�<�����sJ�i��T"���������lwm˚bNK��(eS촂�ʭK��D�z5�n� �8m��Y�N�I�	��B'�����k�G�:��bH狶������VΣ�m:�b/�B�z�L��ݶ䅥�_a��%�A�/=H_���җR�����w<��)��,��j���\�)"ܦynpo�Y���<6���L�FHgrO���w�"u�S0ïj-��0�ƺ�4O(���M���$s/�eZ��[���'�n�ƅ�l��T�+U��: �YܾM�Ҹ�BX[+z�H�f����__�Z|qȼ��Z|�~I�}�It9�暖�F���v�B?D�e�kTB9����D�b?`�����'�Cf�`!x�C�S1��̠�z�W&1�#;o����^6 ������tGT�8�g��f�Ϫ�}rA��6�%���w}� �����~S��_%"8nF���O'e���V�t�FC�Gc�VD�%Ef�� �q��mgH�f���a����˰����y��T~~}��NV�[X�#�BQ�g�7���zj)��,�@��/��t3�Q}Hg���8-�9��MJ�sG��OŰ�-ߝ&2�=�米=�q�R_�۪O	���Oݞ�q��s�����yv���C1����z�zѡ�%��jRfXY	&���^�*/)h�
N�+�[In>��3)n������A�k�N<^*鸨���}�k�K�t.�_�%,�8q^o�0��W�/S?�\��m�c#@n�W�R:��W��j�Y_��aV��9o�9�$�1�G	')[~����L>K@��⧅�y�����۩6��ǊQ�׵�,���m��%�����*VR2�M�+��J��@����Мo�O4�4i��"s0ZCIKQa���sE��ޕ�_h�	�U�H��=T+ۃ��D���p�p�dl�j(�� �.^��|�x����v]�� ��v���W� e5~�2�&�-�&j���ZCO�=��>��5\[����hL���Ħ� �*H�3-=O�c+�^� �Z�
_�������}T�D�遾�W�D�߽��W�[&jWg��|�dp�ux�J2wU�Y,�sQ�udy��Kl�we���4�܀��s��aXzD���\�-��C ��Ŝ?���R5;1��b����Q��;�T�R&� �Xh�A��MչΑ:�I];U@��=T��R��-Ha��<c׌s7=�Jq�F���z�.d-�=�f��@����nU�/+����>n��B��A6�þ�Y��%왺o�^Ɉ���?���W�J$�kї�|�T���,��ycj�[�=�jY�~>�
���X�����s��|���
$/ ���GoM��)�]~ٸ�@ɷĚ��RqK��6�_����ر5���޸��v����*�C!| 1V�X3��;��)g��,k[�g���BeX��� �6q�߾��ޚ"���+�JI��C��_k��7��
��F� �"A��Sb�.9uyOI&�K%kV����m�*���	�^buz~4A$ʊ2z�ҏOO�!0�:1�k�ڹ(��� w�{K�;��:��.��"v��X����+sm�yu;���; �>�@W!	W�޼�����R��4�����z|�Y�v�g��?d0����bRV�G��Y�#S��'���C��'�\8Z7��጗IÔaH%�Z����1��ڳ]`ĥmU�ᝁD���o*�$9	ތ�(9�� ��p�"q��T�2���x��4�y��>��n$��#���i�)��{W�~�N��AK�DR�����45�3�oTp��"����Q��.��?��fCMT���-�e�?<EhlRY[$�y�/��X�8|PQ�e7�miyUR��n�����׸��b���+{�Y��mu�6 ד��`.���IW�8�D���>A�{2���'��Jp�J�A���T�3�$:vW�5���
��2�K��r�

�<ƮG_B���%z��5��Jtp���xt���ġ��$/��1}g�Ď+����Gig�s����L��	J��C��V{�G����}c����dA�2�'�W�#��/�j!�0�㓇S���t�Ք*h��чҸ�z�N�����S˝#3
޿��*,1;a�~f��3����+.��H����X�r�`�L��3���q$���'\�]>G�+ݐڝ�T��Y�&�hՍ�1�vx4�
��l/�_���Qr3�n�H�HL8��G��B����s��eb�O2�RZ�B���C�;��E�ŸH��b�YIRɘ�'i��!aF�\U쒃Oc�mE?[�3BrM^�kx�׉�4����k�t��;��\�Q��g�_=� �r�^jD�b��P:f��RE*Ɋ�w?ޮ�ƉdȤ��Ʉ�D�8s8q�D�U��x�un+��7Է�#tX�����$wת˧����lj8���Z�P1�nl;ig�N[g��u���4��P��ţD��HS2�,M������9��<C�KCH�Q��͞�b͹�&����N��^R5�ݎ(��2��n��%�{}%�V�����d�+��k<p�[�Ί�v����.�A�zG�̬P��;�8��o*a�)�n�!$��ĩ��m�fr��v��
1�ؕ��x�i�Up|�d���)�kJ	�o���p����9v��������3oZ�T�\qx��X�yi �2�Qj�B�ZV�V,<z���#@X<��)���D��LM��ڲ��;,1Ӈ}��^��2,��n{�D��	��xm�ώd�5	����y��g� �F�qZh�E����Aa&�\����+��f��,(��Q4�*��Q�5w���|-�xka�QR��?��\�RK��b}^�܀� eN����}Z@Q���nͷkveptcڀ�'t'����{�<�9��Xn�S�.Z|��N��1�_F�R4@��\=�_�Т�\�u}\�7 ��7���/#xm���7/ܰ���`�����A#��Ulxr	gz��;ZHUN����ɺ�����[���<�d���/1���ވA�F~J�`M�/�]�\1�HҬ�O�#����P��mI!ǹ\�5�NT�	��q
V.�1�4��!m���!�+Tv.\2�P�5�t���5ƺV���4x �l��䔿�'QNuӣ�� �ł��\8�΀*R�*�B���o�7��sop�J��3J�݂2�}�ҷ��谫�U�ђ��`e/Y�`��D�$n\�r�VJ�Tk��Q?fC�$�;�욆T7�+��1�ªd�D�v����rޑǂ�����E�N��Ζ���cu���l`��<���D��B�5Ϥ�潕�&}���-�ܫ�0���D�]u��/\�-�����%|Lm@��,|�(���>{m^Â}��H?%y@j���a0EjX^�C>�0�C	��rd,R!.�
Y3�����W�U�
��~~��=`!�\1Z�I�f�G���'y�Dl	����=kZeF��b���5_xr�#�����F�)+5���M��W����y�gg����c�&LF�|����*���#�y�b�"��@��TF&9Q�J�-ͩ8/��A�S�,����NJ�����%y��M��c�[��'.m��f����-MDV�7e��{Ѿ��a��&�j|l0�R�l�IUS5�.�k������$q��<I����p$~�YS V���0�����Da���ί�|ȟ��+w��:�$u�`���ʖ�w#�y�Z	0��h�p�n6�܍L�c��5�o���Y���lW46�A��N?�=3RaN� ;9��up�3ZىEL�K<�lah�k�H }�7���(W��w_�J�.1��l��8?�d?vV��*F=t&s0?����A�Â�v�Z�xX�E_�B& P2/2�r2���t�
�[���?l�\w:H�j�U7��L&�H{�������$���Ks��g��ļpv�#�4�5C�)|��	L��N\�l
���`Z��x&}�u�Hr�h���/4⩗����uh�M�m��%�'>�yn�؆_dT��yp//i/,�����m�"`�j�m`R�k���A���r���"��_�{%�~s�f�nTL�UvZU�~j���i�J0V��34��$�2"��c@P&{�Y���+1#XS�59�-���J8(��NRn?ww������u�d�"�]�B��E'�kuľ��6|�����Jp��aņ�'���D��k�_�VF���_!��"�|�!�Xi|��v�����?����8���:�����ڥ��͙6�d���\���ְ狛��h�-�s+m��$O���'������{��� �dS]��p��*�`�s6���]TY_	��~�OP���`ڕ����L���X��~�bN;yJ�|l�C*�EUD��1j��9�P�T���XĶv�D���eH����ݴ
����:�Qc߈^Q���
��K�m���/�.����f��/`8��\F���.-�l����)$+��c���/ѳ��^�	�F�gW2�K5-���>ధJ9HG�����X�ږJ��'6�C�*0�::�Z0 �����8˻G!0��2�q��A���8@��dTk�ؕ_8e�w
p���A��@���q$�`�3�f`s}�f��Q'�f�&S�0�I��ɥ8Z��`]���*M�N�1I��$*QJ�t�38V�8���IЭ`a[�d�:�|�A�Z[�$�i_R�}7� <�$2�x�-�/㪝n-��y���Oc���U}�,I�܉�j�F�.(��ѷ�+���L��f�6X�9����D%��k�Kb���j[/ ��lX"��;�ؤPiO�-Vst��LX^R��Z�oBKr�aT"�� E"b�1��u�G�Z��ܖ�|7�'_(X)��y�\���r�i�����&;����=���u�$�Y]���.��vW�I|�
�T�7%rE#���^N]X'4����=�{.@�A�dB�K���,�:����*�zz�aGA�,x���Y��.e���m/YX�"�����!�`��U+�\��J�!�k��a��(���ȏ1{x��W��k�N:��^�-�I!�3C�nҲ���"�������xk���Um�朦�*t��-a�P�cvr)���l<���κJ������xY�{�Y�*��S9&Q>)ƭ*/i?��*���������b�Dk��?���ۼ����z�����l�;R~WO�ѫ�60V��G�vzS�kU���@�H��02O��ĩhK��b�}��3P&A}���[  �.�C�*��DHmZ6k���1�S"U�y�b�T��\A&\g��w	y���ܗ�-{���y�NJP^�2S 	�+`�"F:[� N1sL'�����(��,�X�G*R��a�zs}M�*#C�+�!]±�\�A8bĞ 4T�mE�GOl9z9�A9D�.Zٗ���e��L%B`�9�ߩ��e�X���c��К�	��P�]:��r���@�qr s�T�kXV������������ ��G�'U�0��a�7�!�\!0�O��4ꎇ�Xȹݡ@0�W�OP&�My5���u�U�0� ^��-���
��KNM�Q�z*�?ڀ��6�V���B�s���d����$3���@_N��#U%��1=ه�	���� ��.��C�T��7f���K���8�>����|w�'�3����.�i�Ωq���1�ql;L�J�g3y��ȘV�07]��.<���	���"h�8.M��^>Y���=����kaۢR��<�x6]��EM|A�xK���$;���ƹ������"����!Y,a-�~����rY4�VŁ��l��zaf���������R3H!��l�G�>Ds
>����HL�,K��Hu��o�~؉�5��4O���V���j���+��سqs�� ����ب�@��H�&r������5�TQ	Хz+Ŗ4�Z�!`��VH�TM��Y#�X���)������$�b>4�Yj1ZYtg�IE�qև�`f+��7 � ���_ҥZ��A��e!�'�!�h���zP��-UL��3e?�?k�r��Sr�vt���@ȣ�����pB�5��i
s���m;BѦ����)��2q�Ӫ���֞o؏�,��&Z���F��ܩ0����wr!�G݄K����}v�������
� �P+�6�Hҹ�'aLHؤ�w2 �u����m�<�Ϥ�\�-bt(�Z�:s_x!a�̹�������_����3�x�j1��7v���:�\�P�æB\�!�Lx9�t�5��h���mΑI�({�8��tf@���5�he.ܳM�j��U�3�����ùb|*$�|� �ʃ��c������Y��kD!�aO,�wKK�\��o�wmev��M�G�秛"��lW�D�T 0�}�:���t��eE�-Z(�g�y��q�{�c�<��v'-�榍Y�����e܁hg'����07��z�_��r|���
;ʥ�R?	z��������&<b;����4�9��=�Wk�����|ٷ�2C�X���C1<��L���>�H�%.��^`���J�n�Je����[��B�����i25⡰+6�D�4 &���&�V=�*,�C��tqH���1��y����{<!�!��
��J}��04�4ol�
>7`'Jw������=�5ϲ�k���WI�Hd�}'ӣ��I��W�򘫋 �p���{��t듆���]��\K�8��/w��I4~���r��E�p��O#�i���y1��4�2�=����+l����8�����r��g��3'�Rq�g�]��Qjݴ���D�G/����y��R�$Rl:�7�O��.(2�߶�p����i��C��T۠V��`���ط�'�gF z�*3�~�H1���)��"jv6Irgt����1��/��
�f�݂e���žx� �wo�C4J�v�n��Қ�3ʗ�i�a�D���0t«Χ8|�EDљ�o�v�Þ�T�^�z�a��ꩋ����<"/C2&�M=��0技c�����vy���xU�t�GW0��`�'c�
��No\���b�9�%!ZQS0����Y~�궉AT�ƇL��A�Z
#����s�-wL����X<��6n�Y|�m�Sl�����cj.ɋ���,�~$jqk���`��E[B)=��s���;z��ഴ���!&r��NYp�yF�Y��En]+�i��t=���9�����13$�]}V�}��b�]��|�x
y�H�1�����ֶyޯ4Z劲�v���4�X��������=��+���1� 1��껴���=��N�ޑz��/K�_�ݣAv��]qtJ�0�Gפ�%�z8X�DU�N7x�[y2�xy��#"zP��$��Q����R��Yp��`|(�3����з�������=�ut�^�ڍ� l��x�G��5��!0�I�����R��T��м�ź�J��6$�x	Z���8:!��81�6l�/����5+P?� [�k��?b}��h��k�-�ܵ~��]d�]h�^f{%����)�9�� b3�SDo͸�L.�Õ�2!W����X�FC���`�'�[)����t;�ty25Ku,��"�""����So��i �n�mN'�)1<����rht�%�g>	ێ� �ۆ��)��$� ������:�cγݤ�1�;
͵m��&�|����X8�ϥ���Bݫ�)؇��� t|�[��%��F�6�>�јdf$):��vs�);��`��^E�--�����<�E���J/w���OYM{a��J�=�-&Ǌ�Sr�"��EǱ� �>�ks8ǈ�^P+�i~�x�O�]����� 6��2��l#)�q��f´�ɑ��ԯ�ZoΗ�ǿ�k���ṚH��L���]�%6�[#��L��S���ɖ�w�J�Gp��$UOdl�����W�M���Q���fC_q��Ec��<Q)i(�����KKn�0�+�z�y��S>s��^&#-���H�5]��#�1�=x����(UDl����NN�h@�k^HL��Z�dfoQ�,®Ʃ~	�&��z�S�(�,V��8Y�:�'}Lxx� �6���Tw�[�����P�bXS�Ӈףj�>����Ӿ���d�4-Ɯ��>=TMٞ;��2��<7G{�7d�^L?>�L�|1x4�x�.�q��Fq�D7%��Y��������S�	�;ҽ�Wfr���P,��}qa&�8{�_%ip�`�/1���C��3g�G�zW�kADe�?ھ�(	_�N���.m�}`yC
gS��j����#�d��qk�$g�[b'�vM��a�B;8jޟ �
-(�l��r]�?���F(㐓|��hP�S֏_��֬����L�\�'l��+$�"CH.�����Hv����GZQ���2-��8ȿxK������z��l4��6�{~1�u�$�O�S���V�gaW;� �Q@�Op�������7]L����e4���58a?ꭹ���"���f*/L� ��S1�5<>��3���(�KL
9����dZf��
5l���"p�Fm��;�5�aoW50p��^�?������b[/]ra��*>�e���M��f*{�`���}��{\�5`۳��74ߐ�	=�3�&���)JڐS��ֿ b��6[��^8�b�� ����~ѹ�Q�?��GWZn�/DL�(${[D���.��ixpt6᯾Tl�	��0#��:N���x(�΢2,5	=�ϩ��� �uVǣ�3D����e�F&0-5��@I!P�m�h�2�'��۹~��"~��E ���u�!�3XsHې�p#E����'6I]�ߵ�k�_j�}�1󘶅�O �	�e�.����k��JS0~~�'���<��b��	�?�E-�cx�t� s��Ok�W��k���?c��^f�A�ɴ	#C[����޶De�^��UF1���}1�>%N��CD8�B�Q"R+c❔�?�E(#��!o\�¦J�(Ӣ���dR�i'։�{\U��PQ�A�hv�rR�@dr��?�n@pb���j<�Z�=��ެ�DLk<�?�ʹ��CD�� rM�I�:a�@��*y�A�9�5koh�^Bݽ�W���REԴHk	� /�+Zĥ%-ZA�]���i�E�rM�l�@}H�dU|cC�f��A�3Ų�]�����N�0���1��:8�
�5����@e��۸�Oq��Q��=$/b>�@��ZǊ��x#>9f��9��<�X:����Y���Z�̔8<_CJڬ^�0��0���i���ː�r��[b~����Je�VG�~�u�̧����D�㯭lش���Є��=ް�N�4��~�A�ȃ��Z�yckǑ�:�TԃŮ��6�w�vy�V��\k�Q����0�@����֐
#�	����[�^g��'�v;�Oy�Z���@^����s����=z�V��ߑv"�-4�K����b3Ͽh. �O�4]�lq�q�X8���ɧ�6����r�?�,��/!�������֯B�:��ȥ6.���7h����>�n���`�5_����V�����ZF��C��*� [SN59 ��J��A���5U��Z؛7�l2ˣ�5+��tz�$�d0yN�C�4'`�[�XMwS�@��(Ŕw�p��TW#�%�5	�GZ�~�=�xT�� `X�t�e{�5H�7e����]�����<&�+Kubcb<͏#Ӑ)���R��Y,E�y|uX7<���B��v]��
g�ڋ϶��l��| m �����o�~��k�Hu�͛�~��~�%�T�\�Ėߢ��0��H�)�!M�b��)`��&���%M�x��AuA��#
�xG���>L2���<EEqj�xXqe_B9K�B��&�
Dƿ(0�t.��h�バ"����ʭ6��~#Q�ä�롪7Wk\��� �ei��h�CX�O貼b���j�C��N���Q��g�܇hH6�C1���kt�!��큽��2�aÁ��3�gnV�(0úXLd���k&��Sߕ�{N��������f:��](�%y1kӈ�0��/5�tx��iŃ����
׼J� ��諹�M���Y9XY�q�4�9=X�¤��r5�y�J��:�E�����L�%�K�XQ҆�Vvڙ��;� _�̦5ç���P,�t�����)Ui9)�DSU��
���j���'��q����Jx�~5��=�����*2�E!�L���̅}����O%PM�Է:�J����B�!o��Ԑ����,����L&4��H�h�@���A揙� _W|�4�>ʞ΋15��%E��zͷC���q��3�;���'�n� Ȉ�|3@��\R��YG4Sz)�휝ex*��ܬ��Z"�Z���y����bŦ�&�7��:��
BhJ���^��<o�� JoC`E6�!8�{�S�� �ӷ"c��5/! }]p�u�}���*���s���-��.�6�[9�g6<I16�V����p�͝�h��ܠ�Z���֊׍P�?����.Z��E�`����Y�Ĉr i�U"�~Ƅ�!�����؊.��{(���.07Q�y��ݸ�N�۽������`L�=��5b�F��}�M{O���W�;��$�]��Q�bWEj��/'�ʅ�(�g{�=r��'��yڟ��^hIh��9y�.?`����c5�j.O5/��Eޯ�t�E7�8aM�.�8Ə��/ �����oq�j?�% 쮸4v��0��!DM<��M�)l
+z�t>~x���v-?I�3���Q���}G+��v��a�e��8O6�McuBXp�o�*~9��C��Lqe��z��`�n��Ah��O������Cn�C5�8�@c�&#�A��6�N(c�8k�Xuϔ�!pfڕ��G��Vɓ����}��yE���a: R{�x�-��TX���;���C�-G{ټ�@����x٧&aP��@�M�^�u��c��c��9���y�;�]ڡ{_9g6�_q�J��]�]�V�3�0�U'b���~6r���g�3�$�a���q�@� E��c3�&W��������,���-*��aVY���<o��5��)�������z@\ƣSH�3��&U
�2hoCA�̱`��*�(�왜Hz�[����Is�8u�N��^���T��Jv�ϣ(��&�)�_L�w���.$|јe|M�� �X>zsU�~����8�z�,��{X/e[臶�Ex��UI��4G-�3]�����"��Ck�\)`8�u)�֘g�.P��u]?⳧"�����>ت���g�(�q�K��ץȁ��e(Y�)�w����w���B��K_���� wƹ�	��r��wY��l�R����SfJ���S���i��t� /;����>DS��<~�����t
�
�9B���QIs�q���͞	S������+U�ǳ��"#�2"��3,ܜ�ÞU�Wk�'�sտǂi��8p[�c�k�n�="a}��?ت�����O�`�䂽� �=f.��8��c�.������@"�%{� �ͫ7BS8x�/�r��(�d#>�+�j�������`j���8���5��!�CP�Z1qH�}.�M��AΪ���u9ҩuG�6�F��TO�0Xͯ$��x�Ѡ_6C���w.�4uE�ߥ�X�`���[�b��6��R~���_��/s�j��,���2�Q���KC����e�R���=��q�R����\�~ᡕ��Q��#3��	9F")�r0{f�	�����x T��W�Iq�6���o��d�����U�l��A&�L��o)�J�C2�-�~/`Z�*��[��0�M	ɲ"����:7�f1�w�@�]'�Jzn�֎F���!��<9P�C����jub�@)�;�${}���^�u+5�r=�����K��
�"$F9Rh?h	 嚳R6ģp痼���<�:jCSȾ����i�h�����(�ӎ�u��0��{� �S�Ͻ�K%��W)����A���U���nor|�Q�Y��hRँ���~�ǔ��i�9]>�/Ǎ�~����b�f���릧�0l���^@5��|2�ͅxQ������R���_e
����hg/8,��@��z)���=��o2JU韣�\u��4^;�W� M��ߣ�L��
n:2��N����qht>�c	���NO���04-���0x�fWƢ;���_K�� J��a���Q�j~�!�Ö<WR������M�ʒ���g�������wL��*�������jǷ%3 0�Bq	򕨷��g���X���+z��ԍ�IV�u�.�C-��F��"����Q���~8
l�S���ɏ��ڣ(���W��%m[�Z�`�A���_ZT~�6ܽF��cِ���}�l<0�9�e�r��{�#�����#Ҫ,V`]�Kt�`(���Y����K-PaFȺl��YM9��CgQ�2.b�ʏr��P��Y����y!�Z��8���d¬S�U��/_��%h�Z����y϶`�z����
.�󈬙������9gK��Qb�� @ɾ(��Gz&��]����U/IE�7�����5���=\�ǀ�|d%���*+�%;��53aӊ.|�z���$��z"�K��q���e�}��m�r��5L���W/X���SZ���Qz]��w/J��;�V/��F�Z���(2S�� �8:����F[\�!D8��j`u�S��b?o)��})����z��q�P~�LHj��U '̏]��\{�y�]�B:	�g�>`Qa?VmPʉۄ9Ɏ%{X8$�ۡ����{Q�G��:d0H��x(�["�
����w��a���phW�lQtE�XүN���N��$C���״��:+���K��aI�nώ?S�r%B׌Yl��k�iCl.&�W��f�ydٍ�Q;��n|h�㕉&?�g�>��RatP���Ʋ���������5">�����94>]O���jr�z�Ve(�,~7n��R7�ƚW5X1{	�����p�2&T����#8��u�ڻ^(�Q�J�~��)�D��,;��>��������>�8��O������V5VT�VC�RVU��x�Sm�X��>�S0�������*�us�B��lA~>ճ�m���P�l���F�~��� �+ɫ��gSɪy^N'w��u�,cD��>�*X�����<*���ٸH�Ҭס��#� �E9y���.b�*�d���JhCH��a똷FY¤Z�Ьԑ$�-$7f����f�ƻ<|��br��(i��_�pi�+��ٽN\���m�L���R�e�3���)���C̕Z/y��&`���$�9���O;��JL_v��b��e�3��߶���o\kVya��o�1|F��U*oU�}}�YB���$;P�!c��O1��z�e����BW�Wv�V��;�p1&�J�=И��|�YG��K�(�B8��x@(_.%���P��=@.�1l�]���/X&X�0�y���`���L#�ѥ��-��2~q��w5]`��x�W��_�N_>w�,m{�{��y G�$�?�������v+��#]ю��)}�8�]>"}�*(�OC���$�;���f���k�y�Uކ���c��(��ƈ�bxo0ƅ�`k�*�`����,�|�� s]w���Uf�G�~�s�x|�&�n%�Zl�Z�w�:+p?�_N2U������n�,=��	�5_��̆������aH>��pk��A������|��䁐�߭O*Gn�A���T�^��E��tq�ٻt ����u[����*\��(�������W=����P� ���l6+�B�C�S`01M@N��=Ӆ�y��[���n��/Z<�Ur�#BJ�	�>
�Fw8��k�%Hu՘�±'��8�@��:�����E��L�L*������}�G;pX��*o�t.����>�qx�|���ړh��<�Z�Hbu' N�?7�b��I\��G?w�/�X�>Z��Jua��}V�C����)A_:�N�hbp���Re"�\�١>��B�Y%���%l(yN=�q�9��u����$��?)�d��2e/M+�Ȭ��1wP�0S� k�0-���~c��Y�0x��K�x����O8�{g���N�z~�#��NH;� �<ȹ�,���/�P�\U�,�4�G��o
H��y�,��Y�m�#oI{n��A�	�9[�lv5N~�"B��b�!G�։c���B�0j����ܳ�k(��N(ff�<ٕ�#�^��A��4o����T����S��(�����0HXU�F�S�]Drp��͑N��.��L����M�T^S+���ʯ���i0�b�����y�S���F�c�M}��a�D�)M�e����LmWf�[�2~ӯ)'Z�W�Ʋx$C���$ۊ�]�!�sk��(��!P%Ro��+r�_�������`�S���Z�E[�4VR�C9���Ҥ�x��t�.a�W��g" �潇���R$[0Ѧ��;Ȃ��6X��0��<�I���Mek;nk]z�2�X6XW�`4�t�q��e�����u�6N�'�O ^�@�m}�={F�,��e���l�H�,�H ��/��#j��5b���#��[;�]&���*d��L}v��{f�����2`6��n��EG�����	�gs�Y��

T?"ѡ���H*,%a,|���h�-_��yĜ(�QF=�(4{��*Mj�k�2�W��(�j!.E��p�8��;\v[>&ŕ�bX�Ʃ�b������%�2�]B} {�(֝������K��ܕwm(A�ISDu#���S��SP��U^SC��U�|~ĉ�Ƣ��Lř��엺�o��y@?P��2��ԡS��)mY���8���
2�����Z�������N!�H�Ey��Kz�����b�>���.5��Yʼ�m
��v�5������ �*��ïq���$b�쒧]%7�w��/���zҩY���[��{؅;SZ��^�c�R򆑂d"ͮy;t����k�٧�)?#�v�q���˵���?ن��	�}��p�;�R7oDq/�}	�׫5	�u�s�W�%G�c]'GtPep���8F�I���ەC�`#��+���ouH��ܴ���)��\%� ���,*��\'�\:�Ol���~�ƽ���۱)ꃂ���������w��j\(��%�~'�����Ұ-s)�;�������G���oh+��)�j�Tm0{(+P����R 01\Hu+��"���dyջg�_'G��K�w��L ��H��O��:Q�q%���)���r�.�\��q�7	��c�� "g;`��#�&����ťn��U�
lL�,�_Qh���5�S������f�_ؓ�U!��S��$����f�b3P$��|�a�v����	���{�!�?��#����ԱZ�I�w�#S)�)���
0,�N K|6��h|gk�g���<�v�������QL��%�����A�gM]�Zu,��^�8�����_'�Mm�9
L��ll���^>�3,/'�m���VJ�������M��"��^�k�*'3٨����]����7H�9['��&��^}��GO���WAvv�e<�Rz]YD��=p1S��=�|�����5��]��<�`���3[}�qЈ���3���זD���@s����=������\�>`y��̜�_��K��=�p��#��@6!D���9d���PuT�O�.-��7ghhw�W�>��KJ7̓���Ќu��i��QK��@Ì�S@?��`r��- aD�=��)��*��i�ժ&)��> �w����T �򒰜��;�Fs,��'�u�D� ��7�� �����v����wŚ�SW!�6ñ&?�aت�&qlQ�̽vV������o��ev�f���}�l�!��޿�����D[OQ�8A���ظe���g0`����P��<��j����pU�������QXX�M����h>�q��TX�L�1J2D߸[WD�P��Mc���;�b�2&n�/��E�@ŅM�v�}v��b;K�<6 �i�%ں�c���������~��Z�m�J�I6�7�ytT4��:bto�i����s�+�cR۩U�t��MV׶D�!y�m1��k�T@la��~h ��I���� .+�L�'U��6!_���
�j�[@g�@�(Tr�9��C���D&�T-p�#h�����b�!���[l�f/c�Ѐ{���ࠩfe9���Uͻ0K.I<L�@D�������Jˁ�	�q
���$ic�|2��s��V������w�-���+�٤=�;xx[���S?���=�@����1|��������xP:���)RC[�T%<	{Y5��.C����Ko���їd ��2�ԄA�����[If
� �k"��]_��+#����I��(��ܤ�����|����zَ���f{:��
�o0��J����I#(N��:z�Rx�n�CE���]We������<�~c���-�>!�,��e���w��6�Ս��"d'!�VB����%_�%mH�F��9n�<��o"����Yu��-灿���W?%g��0.�����f�޼P��O�5����h�T�N�|%���Ԟߥ
 n��$��CިRu����9ڦM��o F��;�%��m�~�9�V� I'�m�n��.�x)�T���O��٤|C\	A�B�qg�<C&v*�͸�'?^�|����IM� \�.�KWW�:���n;M``c[	�\�pX/L�78`���:=D�'m��^���>zVV��������|�E7aX�T���$t*���%tp��-�$`u��α-9�
��3��P�ph!��xD�<z�����Y��H��p�ϔ0�O�>6�snӶ��o(�w=����4���{	���
�Q�ט�S'%���s�`��!:�u���~@����Bs�y|�z�S�||�xl^��kس�0Iÿ9��rDd3*�`�ZJ0\m�C����<R��y3�4|C3������f�9�$��xl�Xط'���p}�'�A�'zͿ������^�wq����+̶�ꉍ'HY[z}�
`��?�1#��@5"C��xt�3�l��w�ދ����@��s�C`�}��)��M�z��pq���������Z�E(ܡ��@�������*o���&��꼗ہ�f���_�����(�,ɽ�=c>�=i*��i�
;&{�����?�\�
ĸ%�����'�5��'����3d�W��h�1"����0��Z� j�@�o���2z�3O�<�5׀�
�$����kW<g��xɄ����102��R�����>��<S�;�����~�i�߫��?}#+�*`✺KM c�������|f�'� ��>2h��@�R��C8������l�'�.?��S��0�!�BR�����Z�4@��
�j��C?;���ՃY�wC��o� y���C,�,�37������n�@I���A�q|vi+���&x�6W�5������"��~K�eq��Y��G|gB9S��4:��|�@? ��L/���5p�����D�u�3yg���<u�5Z��7��S_��9���ms����) �J���g����Pc0o����T���?h���;��F�f�X����hXH|�B���"�m���d3z�vq t�]a,�>�+�+�Mt-V�H(���}����扛��UM2DE�m6�U��3򮢫P
D�y�9�XfAo@������sہdD	��Ck�a��
[���$$���IM�p)/�-B"K�dJ��Q�������夘v��t�v�R�E�X�K����wP��<��}�թE��7S��t�V�2Z�����=C��y���/k�
à�O��i�/a�^MѪ�ߛH�)
���c̉͟��Oi�1E\�T��K:�⬈���A�P��>,�D~҃�*I�g<B� �R���:�d�Kl�Ɇ�[tt�B�\d�z��p�ٌG#Q�u3F�=�*��	΋�U���w�?���r�ޣ�ZBn��z���\v�������}Ҧ�0��Q�d�����bZi[eL�Mw�T@r\�G�YR�KAq�Cc��:rG�`��7�p�VP[�R������@>��#>�\�CaZ�́�fDWet�T��:��_wj&�|���[r[].΅������,(���jA^� �����TIc��a�����AZ'O��!vdC�UM�;�L��P�}�}��ĕ)5��$5�J�T�g��a}��1:�+IHNƢY��:4��D�o�:�2��u����>��b&�H7���RY
8���Re7��O�K;�����5,A�|�X��S+j*�L"���jF
����3�6�@6��Dљ*��l�^�֢��ѫ\��@��`�)��IW}
j��{��sq=?!b�I˪c$@�+$�:^�5��8�(�F��l��E���� ���I�f����IQٞr�F�dOB�:Z����M-#�Xe�>Ŀa��#�L�C�6���Ň�ͭ@�/�ܳ6$Pu�#N3 ��ַ\�!�}������IAQ���Q�q�.���*l��I��۹�R�����*��\��J�ܭ�iڲ`�o���7��!��4+�єN"n�W�\#-6�ƤL6�M�x�i��+�z�`�TOy�&:�gN�@Ĥ��c��`�ȉ摹��[,5_Pw?hvU!��8���]����5a1�(.��A������FCif (6�� ��Χs{#jS��+��
�;�Ϭ�.�S�&f�m� �[���VV?�+C�9{ʡ~�g<�I|���-#� �v�f�7���>�T�L�6�F��ո������[^��|Bn�w���`��t�v�w�j� ��6�������e�c��C�G:�a�.�.PU�;��_�IN9�!#ע��jp���n/:���}�7�a*���JN_��l ��J:�I�5鷘�J�5u���c�5�{�Ǜ�$�<eR\l�M`vϚ`�S���e���b�=i��2P�Ub�Ӕ;���n���
��^y<���)�R*��i��7��N�T���lC���rG�q�lE��j ���J�b��7��$�_'�iP�/�9Y�_����2�N�f��.����.�z1��z"����%�����p5�T�)�Ћ��j���fTO&Qd��G_��������H��n�i ˢ�͏[a�C��2�T�3<�\'�Z�aGA1�'I]v=�P~���?��[�T����=��y��8�z�[~J�DN�j)Q�&�TB����.[����t�x���,2]��{�C��>9u�5� =��FnW��;2�3��P[-��ϝMͥ� ���
,]��q����uT�$Vs��`�K�k�y��c���T��k}�4
�ݰ��������$}#�©U7�v����H{���k]+*w�&�hb�=�wpW�����S�^�y����Otv�HS�ڥ���Eu�s�Pi�|D�y�N�haK�t�RT�;O��D��o���p���h�(�\;:�q���w�&�KW�cn�^ү�l~�=b��Jč%�wo��4��Wu�'.��_x[��������J#�jK�S�<(Z*o�ٕ�X�z@�'�9�vgh�g�IS�(vэ��)<
o{&�pK[���,Q��8�S)�m��Ka
c�*��e�� oeh�.�6P>=C|�5-������m�jM�������7T+=���io��A��e++���ZS��ek�_bM=Y�T�#�D�FJ�M�l��"���q<��^�4���#_�� �R�W��*�o	j�����2��T�:==��Z�;���Ya�H�N�Hc�l^f`�651X�vT�Y�����	T���ԛ�Eo.�/��ν��?'B�g2�i��H�D_t�"��2BF��|�璉�����G���o8Qˠ��/��2�Y�Vsg��}��㑜��')	�=��	�J�������w����ʡ�,yڻ�tD�/V!4&�����T8.sU�ɥ�
^
����@:�%�{L�S�=��,�Wڻ���Q���,<���I�O��p� �]�p7������%����0���p%��"#_��߃�5~���u���	�4��aLK��Hч6� �+9���L��hk����I.����_�r�4�S���3"�a�J��B�z)�9�O��a}���fu�!�Ő~�m|#&�,���'�yӺ�>���}�ꁴ����5TEC�D�5ھ�{��(���A�����f^G:*Y�mv�\N�4P������V?Xζ����!v�+I��k��?Mf�k=���T������FGq�=-c�Sn��6Ԛ^?|����t��D��l+�B^������f�,�+��P�[� E���*���!�-�{��@� u�v���J�6/�R��5ǪX�y� p���4��%Sp:0+Q</.�/X�}�JUU���=��kb�f3>�&�u4-R���;[�F�,�D��$h��$��#}�G^r�-�\	�eʹK���x�=���J�"����x#��cҠg�s2�9+Up��B/$`E�]���Y��(2�� �"��Mg�� ��q�aS�i~x k�ؚ�CQs�KN��*�'A�n�F	�:���޸�.L���#��h�T�~iXy^O%�8j��<}��䘇P��x�;��
�H�8`ˊ�|pݴ�(U8��n�=n�Y���h� �+s������ᅳ��"5~�$����/s�����^���[��ړ���X��ߦ^���2fZ}�& ���>،T�����.q��`y�
Ԧ�q_���'�4*dɎ9v(~����{��i�E���f�F�u�<%J���$�[�:�֊f׮�vfC�w��5���K��f�����(e��Vԃ�Mv�D�h��߭�*��ݰ��瑍7�O���_{w(�E>�-�$����M���ǜ#d�:#�ϛ�5��T�d�B@�wh�ߑɅU�>Y_>�(HGtV�c���Vi��\�T)8}���P-x(b�e2�lQt������.�E��'Cq�p��3&�e7��!őC;�#�3���:��"��\f�s񤩘1g�z���cħ�{**D�v�P�!2��`�0�.۱Р�xc�t�l7�q-t0j��N$�2�4�՞���
� q�J��
M�x�)ĸj�?�E�{ӱ�6H��2�F�:��8y������{ޑrx���q'�4ĸ��r3@:�-+t�emb���`�Y4ЩP�0��l��Rb^�;�J����@����k�J1M\�	�a��<��h��&^��5��d����Ų�
���z�,&K����3{W��(�2�fN��$��^Ohf�?�nR��1?�8 ���O�R���E��TP�a_��ND�!x���PPn����;;$�h=�zQ4��d�{��8�֜Ika˧��z$�ǝ�'�B��n�S��G6V/U�D���Н��4$,V��N�>k&�C�XW��	N���ܢ�(!ܿ��s��$Q��5��[�#��dްs�,��3�I1���I3��m�m��O����w3���F�ki�W��̿;U�@A�����"�6�D�Z3����l�_�P���b�Ex/�P�kʘ<�8������E�qn�����|b}��d7���3���*�rM8��dj�{�kȾ'z��vu���v��ķ�\�sw�mH0@W�vYK�*o
Ǆ�3���Mp-�Nr�Δ��o�-�2xue�el�U�D��%���.�Owy&��br�J�N�O[a�� ����[fh��ݙ=�B�cp�r�_:�a��6����޽��H��:_��8R�����LX��p�΢�{Ǟ;0֬�Diҕ�L�[7�o�V�֨Ӗ�y��f�9�,�e @�)�Z_�C%�G�S�O�l�vE��Hʐ����`s̄:͍O�:�ZY�{-A�	�T��Ԛj��Q�ZY�ǋ��uGԛ�ic`,\�^���&,�6�)j�f9v*г�1 �V�V>J�+ҥ�ўTܰ�[�bΡ9V$m��	��
����T�����3���=pd&������`��h�nL��+�)t�IJ��P�'D��[����,J/��U�z<�t����,����P�:��UO��K>l��>�4��e?�f<��9��geU��fA�>�����c�E�&�t�N��L ��W�8;��_��&���H$n
'0鶭��J�τ%p��F7�20�i�r+��ΡvO;Ao1D�>C�h��~9�8�����6�jS����OV���[h��z�cN&"�%�y��R���>�zl ���<(��z��=N�u4���M��kQ��8��P>�����{DD~�1`�H)�d�O9#��9�U���O��H_y�����f㜕q��2M��Ɛ�Fh6�`��\�x�o1���L1�rO�C
VL=���֦�h���E#2����k=���S	D�	��D��p�$i@�>����h�d�6Dt��~��l n+uu�Fϓ{W��,�Ї�,&Q5۲�p��Z���sא���17c~�E1�7���˯�땣��je�V��Ƶ�S��V�xZZ\���$�3�{��r���[���#���|��R�2�uaZ/Ԝz�A�<�XD:ՆE���$�V^��wp�~�:��Z��6`��C�T����3ԉ*l��|�m��K�)���l�G�!iZ b���1�n�^R��0UE���<tD�`�<e�ΐ�
Κ����u!��<X6wP"{���m����K�J���oqe��u
ϼ7,@:i��[�n3���rz`����x�6�Ǝ�HK�U�޻�k-b�A����Q�|�|�����:��n�3��o=����o�͠�bg{[L��gj�[�s�1I5���c��<kn� ̴Z�6�	i��v$�\�J���_��S���G5?�m;�:]l)?�?%6�ɀ(F'�!q�6(���	���C� �/j�9ν��±��Չ�|>ɡyA�^�)bs���(�R�P��.XC9�[��N�F��w��-!?-�wN$�J`��>V��*���s
qa�ځ�,��񳀃ij� �� ���N{E��y�^�Ne���ܯ��oHe��m�4~(R.s,��#HM�����^�|��!��LEIl����d���v�|[�iO_�#E��?����| ����Rt�p�� �O'����5������A�
�J�j�X7^Q���E.�t�:<U�f����zm���c�!9�QL�3�K�S���e���N�f=a_d�z$XR%�h����$8<h���~�~\:��iN�ՀP�����) �����\�,��[���*���EL���^H�����a`>�<�����k��
�iJ��
�_!c[�*�S�����hb�N`1[F�6��vPKV���ju:����� ���:_��ç��Lפ%XК���Fͱ��)щ߬�vuCC;:���JR.�q:b5�Ƅ�#����%y�
)WV�4��L>f�˰���d!o�Ʊ�����X4~�CW���.����P8�=m��r*5��b j������A����L�{��������Iϋ4A�ӌ�/|����
���F�,kz*8�X�B-
)|N0�st%K'�e>��U8'��'i��� �����5���K}�AQB^y+_T �|���"E(͜Hy��q,!r�A_�N)�S�\�x�&�3z��"'[���ob����_t�L[ُ#Y���?���{�`��K���}Rg�«O�m���A��	�_Χ��kʿ��Vb��w�akO98�%R87Jb�*�~H������*�gh}�mg#%P"���,�-���H����Ǘ��a��'��>Q/��-�>wi>�� ;�`* =�)�JVӽǟ�R]f�"�Z� Ps�Sr1���u:a�NL�J�p$46H��Og(*�3�y���똒�AF�K��y(�O�ކ�x��q!ӄ �&�~ϹRyC�{d^��{c|xv0��+.���'E�8Ͼ��@�K J1���waS�%�׹N��ӌ_�i�,4�-!��!������-W�ɞf�hf���q���ߛ��������r�9�RX@����
����j��SL2q=\E �)��_��+���0�$�~{CM{MH�8��)!��҇	I����yP]���f��5��
�3��:j��_�&d���ui\ŗ��e�!.>�ù{|�C�ҳ�M��!�O`�7�a��Vȡ�#������t%O��R��E$x'���/�D�9�l^O7��X�q��T�Bc}�V:�|�RpSp���j��_��u���=q
Q�D�Ql��)&�>٫�����w��j�aF�<C���L��@��l<���2k�E�@�o\Ɖ�hj��w�N.E���g!P�B���,OL�3ӽ̲��l�w�6�B�E,mV{S ���;��![�C�������8^���"�����jZX3-4J�	&kh�p�����7-�UH����k����[u�>Z���jk^�@^�Ryw�7U4k�����E�"��f31H��SnM���!ֺO���^n[�y(�9�2Ji�>?�Y^��	�1/fe�|�<�d�j{�;�c�BZqfEZe-ŕ]M��z���¦?�\}����MZ�*�!� r	hk���;F�'2��E�:����R`�x�SQ2Ɂ��~����@������5����\�����~�]��YXiP,�-��d=�Z��"�w�(f@�J�0Z%8�	�y�諁O
GG��-�]����,w�q���1��=i�Z���0c�&�w]� ��
�Dմ���T 5�J��ѕ2pN�P�"�b�\�d���֩�BwYb��F��dP1�<����{EP��2^CM<��wP�S�;��� �2��G���?]Um�k8�b�?�cj���{b��w/�'!V�� �.�	�U����Gv�%I��m]�,��j�>���F�3�G���H�灄��~�����_��VMBGG�Ī�߱�3NPS��ؾePu���`��Z�٧7̟�d@�xޮj�ÿ�r-��v#��N�/ �krmy�/�B.F�
���G��P3����gG	����,��;���*u��wKUC&����%��Ӊ�Xg�P!���[�����l��<����x�'� �F�V�bK>Q^��_?�	��&#3*����x�ɛx�Y���ސ�����������������LU����#f��}�T���,F۶�`
Ƶ3"m�� ����&�Y��(q h_/����~�m�;���F2�i�	5�;�$��=v�H[���a�1�H�]����T�VN%Aۯz���#P��b$`��C�\G�Q�c�68W_D�c�,k>��|4��b
��sw��X@�7(��gs���l</]^^TIcl�s�OU�\_woњ�©����|^ia��q��o�@�	����Pϛk(�c!C0�n�QV'��q-?R:{Ɋa�����0�D��ʊ������L��I����Z�J�<�1)cW��X�l1sGAIk�{�4��q\�0Ć�o.�Y)�f�Lځ{z��Ő��}
�,5hn���.B���A��S��I*�FG.A�*�@E&�}��69�s@��6^0���E��<nޫ�ǌ[�C��n�֒Hu�Y��:���[:�ǽcb��闧�����+����� D�����v��!�	�
��uݛۆ������2��?6��<D$�>��=��'yo�k�{���BR��\�gR�1�Q���S֑�c�4�u7h�Y�Pڰj�@o8�N_��P��3'��ڞ!3�|�[%�0�����׏Ipc��>�,EW �����ֻNB�q��PQ��i],<P	r�L������x\/9�`����*�mUQȉ;�e��=-����2�M�&�t��ߝ�uQ�Ĺ�s$�D:�3l
v��B���#�Xa"�d���T�)Q�ٳ���m7RUZ"Wf/�,�:nj_��<�`�ze-�س��������(��� �.ߪ�f��T�%�Ar�r����E��h#�-��N~�a�"-�D�i��
��}���6># ɑ��$�8T}UZ��%T!��*�<�������
��䓊�r�,r@^/���5$(�D��TԢ}�	�[��,��� �*@��}��)'�!Ow�a�.wnd8�p���+ۏM�P0�3�
�f��ZҜ��J��fN�����?Y_� s��]�!3��a.���e�-y�y=˛���HXmE���ض�=G���1��8���V��ª�{��g7A!kE�r���:���26r> ���TJ�A�į<M`s�oK�ŋ��'��=��qv���t�j���c��w��ǫ+IG
8�Z���c��O��+Z���A����	��g?Bw��@��6�D���������?����
�X���]��~�þ���]����h**���lp;�	:���W@�j�2�To�[,�������q?FT��,��� A�}�A �Dǩ��0Z�}���8��de�|��(% �X�C����}$�p��Ķ��/��>~ơôN��{q�	�icd,�O�L<ZÖWo=�@��v��tpo���L�Ν_���԰�
��ᡸsݵ��HT���嬃��|�u�>|ݶ��2�;QX[]j��'�~���9(N�����f%K�ED�E�k�-:a|+���\Da�� )�@�Է>w�����T�<�I��
��.���X�����s�zur^��G����5d@�Բ=H.�&z���`'�1�68A�����Q|������P0�.�Y��0AAp��XE� ~(������Q�-O0s��r��x1]X��0�i�\�3 \eoƙ�ϭ9{gp@�>�W����TG��s���#T��	�A�� mN�pTZ��r��>�O�`�j�0g?7�0�Q0�- �<��g�����m�i�H�&�U�W��4m�&��D#᱅%�
�-�z�8B%s	V�{�dg��^{����?�L��,�F1�	�]&:ߴ*�v T�18�������R��v�<@ۧ�rE�JE�P�e�YV]2�pf�r@J�3�uȭg�P1�����]*|��N�РM�Y�������_�xG1��0K�;J*��Q��#�\Å��(3 4��,�d�ŏ>NЇ>?�n�#e.s}WҫsA��ڬ�3P];6�XkB�|�*o��	��:V	/H���B}<xfNu�ʻY�%!� =��ZX5�Q9�N�^_4��2@�if��鉾��i�x�D�e���F�"�|�_î�������#]\��U_��Y4���f�2mU����?�����|(f�����ӗ6�^`$�8K�$�:��G������z׽x����>B���������7�՟��Ub���nyH�.�t�A�V���u5gMӟu"�1B-"i�UD�w\`�W�ҳ#�Y��"F���#}�P1[5K�_L�\NۓE�����<¬�Yw5�}3� !\O�]W�΅����eL��$�hq�y�s#�����O��	Th�B�c(ԝUq*c=�TRR}_�����6N�-��x5���p���`�N5Ǿ� }
����ȴ������â��4��4��5Q�ggۖD��!����Ov���ދL��`ề1l�6�ԛ�av�f�u�W���^`C�-O��4(��T���o�ҥ�,YY-�L=v��r�f:&��w��#��"`��cbC���3:�r�u%
:���'��|�q�&�`�/~���Mg&�d,������v�j�
��$m�E��vX��sb�e�01qvi�r
4��1N�a��1�b��mƊMN��m 7~*ή��Dۮ��o���C��P�6�Jf0ueFv@g��5�5s���>��G(��n]�}�C�PD*e�`6���-��}d#�J�¾aT���5?���@(0*�uE��WYd4\�|����w�*��ӟ�!g՟��9M��z��VD�6cI���K6����:�Iv�;3a�������e%g��6��˚���'�%A�붳2P�́E���6R�V���+`2^�������3��mE�:Lh�ۂ�����*o�N��4���RP,N%O\ˍ�e	�/u�@2��z�jA�7�iHk2��*�������}�o�~�Z�m��.�x��K�2�3R.��G ��wؔ*۰bT3�dWPq�Ti��f�P\#����4�3s��%��<2��ۏߊ�nb%�uǛs�*RH�su}4	p�H�#���G���+h\�L�K3zUY���{�b�M�s	����/��I�z�]{��sA�˝I�}��~��X�F>7�ov��`�e[��:�2u`!�����LLp ������9�Z���.�M	��>�^��X���"`��\C)�KP�X|6L�8_B��>�t�s�w5���\&DS/�g'{�J�.���=t3�k�I���j&�ÕA����z�����
�T�*%벾��g�ț�֬G��0�\�;�6B^s�e4�ʶ��<,�'"/�FA`�;����+P��G81�������N�l;tDl�udZ�iS��3���q��It�T[_5��������\�b1d��E�f�Eau��x��h����vE����uz�L9�v�*o��lt���sQ�SO��?�4�1�)u����X��Y�{��d�/)�������{)ﮮ������_i_ r�Exx��7����o��V�\��^�&K�*�C�B�O�K��ն.Z �����x��^'e����Q��灆��$GuL�Y�zd�W2o(o�ǵ�q��D~��e`����M���BD7��#��Qy8�>b��u�љ���ce���i��\�R!��A5��|�;���[}�k��Z�m1���Qx��ۍ�ip��pE+F�/%('c[���oW�,�٪_}6�Z�ʜ�֢���
���I@��G���c��`
V��Q��6C�tNh��V�-H�V��j�H���<��RM7��x�zJ�w�0�~��f*sg9�Cw�>�<��ї�G�}F�񍇯�:8b�����H���fC���.a��&��J�����ˈ�M�A�'M�3L��Y���]��Rp�]�;kW���
���d&��]�;� j��U�7S^�;�U�|m�R��Dcq
lmLb�b��	���ƌ��S.��`O�a�Ps��.��|]�s���L�5�۷#��O����s�_W���$�܃~�_Dm�[Ч7¢rf�k`j�~	��g6���Z��8��n뉭����~���.�g੩,����qB�M��w�g�n�u��t2�.}_���zƦ9A��]a�P9�D��U�W�R���;�F�q��%��	���.�FI���ܳ��R?��e�|�,	�g��R�g�;�4��#�*��s�/��bcdգt�1��N���zz(ib�lh5�շ5�5�[��L�
�i��	���,s-�l��RR����uv�au���iHL�06 �k"��#���¶Zɻ�.��^(��Qj/^i+J_�\�����ڙ!=��k����v9vPy�uI`݈�A�Ɂ�#q�٭����v��u�0^=�-��=a�Ey�ϼo���kf:�&��N���J����s��օw�ؓKRYӦ{M˸��S`�@�DM$��C�&�1�H�7�w{3Df�����8)��T4؝�=�aoM@��h�V���(��S�/�� �LV`�� �}�x����,x�xn�"��#�}\�vbЩ�o����TFP�S dP��.�'�޶�kY
`���j�u?UA�B���c��&�<��6����a"�Uv����Y��cZ`��E ���x��k�$����ɻ��:���(:Q��q��H���E%Ֆ������!BF�y��Y�$b+j�۶ځ���d8ɀ�0�tn��B#�t;��i�c�8��u���ս�d/��S}pq$�t��Q����x�+N��F�X-�#�m�ʇ����ki��K��Lޖ}m)�
O�e �[#\C�maf����H�:W]O�o��ym-�,�?����y<�b`��-5X��7��_ѬOt�|������\h�
�#>a���:�L�1L��"4������y���Úa*4�bq�a�({?7J��@�����"a�G~�7P���I$�3汈Z)�e�AM�ax�h{��g
�n:Fg�h��:�0_"�w��,�6U��s+o����Iy9��{Ď��Ά-|��p�E�X;�������D�>��ҘS���h�RB��M��Ma���G`�(�%u���X_X��t0�:�4酬�����`��� 0�"�;�X"�R��V�skK�^���%��S����ÿ:�1�{]c8y�l��5'&Y�6�ɸX6z-���]u�H1��������/�U�J�#M�ȫ/��������E-�	<��N!!X�*�l����w�ĦuF�����c$�?�x�~8�q���gVv�&�F��f�ҪwJ-���+̥�P�6[�-v���r�ѯ��aY�J�R@�s_Y��Gn��0HO-�rJ��pV����NdZ��$��SQ @΅;,ec'
 �����<��.����~����U���yJE�Ș>:Ot5I��9�/��y"��&��&���D��kx@�b��rЦ.���.���Z�������Ҁ��J�=��ˮZ�P-�8��M;����34Dp�X"1�]W;sɣ�.!�	��~��/n<��������221���'����I���C*�<a�����F8��*�2ڮ�=�7���8i)խ���û�Ad�V������!����^��v�����qc����J���<�	��WS�/��1��z��݆��Z��&�-^�Ț^�
ϣ9�n�"}Val�֏z��t4bz����3�? r����c�6�=񤱌��	6�H,����gv���{�Xx��(m)�o���ł�\x�;��n�WS�X��/׵�=�'ʐ�"O����Cx~�C_W�������)y~I+Œ��Hw%u�'�<m]����M�ʚ=-�k���&������k$�j̍�'6��te; .Q��J��+�F��n�0�J�U�>�}�kn��m���~�D�p�P8�t���bDǊ^!��2~v�⎴y
�J̾/�V�f�Ŕ4�)W`"u�^=��&�v�C��	"-�5�ٓ9ܟ��z�+��̛��Q�����������tX.���CuroF��c��x�Ώ���	��d�n�]�;�ӾfS�O@� �uAǴ�?(M^����6���L��A
J �mq7�^�,NE�(vL������ �R����&P�	I���Q;��f���P����t\�٫����ŝ���O�ۡ{^�7��RC��>-�o���q_�,������1eʐ�=K����_���)�m�j�Z<AJ���*3�1���{K2�}�#
z�ƻe���@�M޳���&)^zs��H�i2���_�fҬ��K` ,S�D��������9��a��?��bwP[�����Q�fq��_�_�g�m���Zv��L#,���$�20!;��jS^P�П��]?ZP�i��+0sճ�
n]�,����::��x�Jo`rԅ\�A�v�N����=�ٚ @�zfS��
<}�JN���+Z���9��.fT����2�,��;B�8nv!1]��՛P�2�V��m�RH�
���|�埁|k<,C[��{�Ocgٴ�!>��ALX��'��������;�e�I����mv�1�lN(}!ƃ���#[yK�}�U���凧0��;M�4۹�T�t+�|�%e�rzK�vg��� ��ѽ$�l�Kpr�;�J�m�ڇiF3�O��9恌����2�ی}$���4مY�V���Ǆ��q�: C?�JI�D���f�WRU��k���!�T�#Q��U�^��	PN�����B�ib_�m���G�������J���Йl3���0�#| Ш��W�~�����HGzТ�8����b'[m/ϫ�������*c�p�Z&i������9χA��������=���:��6�t���qxÊZ+�Q �N�ω��=������3���a�:��h/voA�%(E6���ҝ�A	W,�]��CwB����xA�c��J{���Z�r��M�;�0�%X��I4��U����^���o�y��l�=�$y
q�y��0����u`�������`%�c�*��^Wyl6+(<�O銊H�:)����!��!X�T<{�,"���-�dA?S]3Q�0��S(�(�T�(�9oP(#�r��pl��+K���jGP��~w��yT+����m*���	_��$9�u&ڞ����p�9��� V�VLe���q�9�`�o��S�c�&D��]'û��Q�h��M���KJj&:��������r�%����C��Y���ݭX����鵞����Q�"�DD�F�g�[�r�6���w�!�t�w�iw(㖵���u���~�;�Vz�"�zy�������.e��:}����A/�A������gy��IH$]��4 ¿ �K#��������I��������f}�̧\'�Ik�4�0f9Zت� c���F�Bяo��Q�r�D�h��Q/��z��>-��_�ܤ_ˑx�2*\X<g�q&�8_ ���`���Gc�6�x���[���ht+�7�~��~��M�{M���:0�v1�*�&}����i��G!4��XX�d]f;�� �>ҧ����pǶ���d��ə+���Rr�P�Fǃ]2�+��\�4;n�}P1��.�=�&�g#��C����"3n�⍄�-B� zM؞�R;r��?Þ�51�0[}�"��~Z^�_�m~?�A�{����}��.��\�dG�`/�P�1���1q�|���O�1���;�X��s�o?}g�ZsnK��!92pN��*���0_ ЯnItgb�����ت6t^���-ځ��]��4�=t�%���U@ ��,���S�|�T7�<�'tz��'��[.����%O��h1r��D�S���%���f����yv����@Աj �`�2g�y��()�7PO��Q�wD�\z�Z�^b~�1���{����:ް	�{�~Q��%sʌ$1��g؂,�}�M7n�� (>�{e+�B�9�V퍩���tW��+8$(:� �T�.������d�b�%1�� �`C 8�e�M�B�-l�6)�_/t6bjXh�^��;�k*��.q�-��[E	�z�:��U�P��A0���=�}�r���򔩺[��~��i�9�e8��^Q�������d��]y�)Ѝ_�2�K�џHf���XG'4��H>�c��~T^�Dz?E�%�nI�^���M�9/�� �;�M�O���nXr=��lRU�p�^٧t�&� ��_5�nP�?��ҏ�����zd��ě��3�m�Ù�(�"��B���:%����XŮT�~��➺�(��:�ݗH�uL[�R~"��{�@�
��z��|��EȞ����!�Z�����mj����#H QC1�ݕ���a0��fo���)SN�b2ӋBm���;�EP/t�K��{��vhg�f�F�j����hR� �{9��v��F+6m���.��/�m��i�u�kir��7���>�(9'݌�*1��cӟM���ge�|Cp�[(�R�'P^��K2�0Ċ,���h� 2��M`XǄ櫌�J_y��T��Wn9i���ɿ��&�Q8�t�A��'H'�Q�"쉆kL�~(P^�V*FG�Ӳ^Խ�tl�zu�lzr��O�������.4�̀�n��l�k�0�Kᢛ���&�����|��;<��S��\�]-���P�N7����WQ����B��\&u�.�~F����t�O+�u�%��Z�e�*��.��8�]p՛�$]�)f�3��s�S�4a��҃2EO0�c�,�vO��+ղr�PN�T��di�rטUrz�R��#�
@�Ї0z��w�q�O�O㈻��.���F�{�õ;B:z���QM�IO��}gqn=�#��c7hJ0�h�V�8���xlHGp���6�/P�|��<'k���Õs16/�Ci�i�Sn��U���,�UDH������6m�u��*M��j�}��0fL#Ώ_7������o=���L�ߥ���<	�M=E�L�&�̘�|	���m8�3&�P���k� �-6�d���/�Q�`�r��s�FĕV�h����w�"d�)��R����M��	�H��Dq/;'Cle(s�L��1��>��;��_*-��LLǆ:����+�}	8q�M/�̣&U�SP+�x�x�
z,�ȝo�Q��Қ=��|��/W�\�8�)��ю.��}}:^��O�۱��������t5�L��0�'��Fk������'Pxs���{�)��h���ر���Q�)��v%���`�����ww|���J�N'�f!y����1��g^������6�R�"A�QF�f��$��I��ֺ��E84�+XK�@���CY|t�p�ī�ej���D����o�H�T�1�_δ�`�|Ӵ��1�C-�$�0������h�I�`�;#_z�J�Kc��7�c3����#�ց~2`	�^6R|W�<�QX`��ܖU8�k�����'r�d�Q��p�R[�����v���qG�#�����n�V2��%��蟋� ���*�E�-����vL�M��TԎ°�.�'-yJ
��F�3��6��k!�`�q��l���@�����d�)�g��w$��_��A���
��;���k#�xܙ[ͭ��L)��"�k�3��m���R� ���*�?����^�B�on��Og3Idi}�b,݉��7�Oui?�6+p�~[�Sz��]�D�.� #ۊ��W���!�o��Pk?�sPj�f#������p��@a�{�gV��U�!�SW�CX�0"A�V�[��T8���˘S�ǭ�Y��q�1��c?-D��C=����:����O�O���l���D�kU�ʢk�Қ�ǣi�4����2x��Qn�C��K+@�5��g�aR@���i����V�y;8�p6�y��Mx��!k6-�`��ӿ�S�?Uv��D��A݉ �����Aׁ�k�� `��}VL1������G�A�V�%�]k��?���5�G����QF����S���9��)��L_s�6T�<��Nw"cG����<i���G1�k~�)�6��H+����� ��8^�2����k{"3�2�j��CNY�Qy�����fE�?��A�~#�$��z���k���PZ;�97�m�QO�OD1�q�j���:�G;-pS�-,�����w�w�8&"��dAy���h�V/ИU�H.�ڐ����r�<k%��T#|�>�fcH݉bo_�Ѹ���%���w�s,4�,n,�V7`�x���Kg�O�jYO��Ƨ�*۰._��b;�.��m2�=:�h�7�i%*��!s�D������V��TJ:f�}�C�������A���T:��r��(�Ԋ$#�J)��-�����]���j7Bvj�=\�`�=��(y+un4��&�o$��-G�Q����"�+�IO(P��56�d���}��o����V�n� ľ�
V�x���pp�C�p�})۬(��m���;���܇pvF����
��t����x��s�;L�疦DP귄�����y�c�Ѻ�HHOk6��ͣ�o�A�QA�޸M��:��/��f�'y�''��ͦ\3��4�nW �qገ =��X��	��o���1�ݮ3eon��*��Pjx��io���M�&O/>߱b�>P�O��t8
'�{ېC9�;d�o���͆pGMe���᜼))�ҧ�06T_.��Z|�ʹb{���TAqW(Q��(��	K�c�9i�(����׸�9���H������(�;����Q�ߵ����=����s���� e�ڟ2s(V#f>$d��%�c�# K�u�H��gB�r�"�2�����Ҍ���8V.�����~��됂D�Wk���J�ܷ���0���[��p����S�x���(�K�
�����˜} �+����wT�Y#�o7-0ˍ4{�uy0Bw��ws��u��qc���� �a5���T	A�$�`%m��OeA�3Ѫ�@y�kH8�����v�oÏ��5m��Jm��� ��3�j*�Ġz��<�kPx����ɭ5Q�|�}�Y��.E��jɔ�	�fT�j�j�T�7�"a�!�$�0�Te>����⊬莣�/�E�{
Ƅp�G��@q冢b��"C�`�83~m�~�A���nr���
�@KYq�B��Uք��z���>�r߆u�;��a�ͯw}�ɟa&Z��Ԩ�>��;e�["O!RO��2��v���O�y�)��/�v]\N�{j��1�谳��$RK^T+��^ӖĪ2�2U��}lH^�k��q��������o
tȠ+�ԙ}>zh��"�����ĺ�J�`�0eI�
GW�j��V$h�_������_�+��7���8j�!�O�vJ��뱬&U�W�V��	b�z|+�E�.��"<\f9�J��s(�O�83@3��% '�\�E쏈�
�|��4߄��O�A}�卂�S�
R0cs�˭��
���L�h2��D�ƣ~s�'_�,���"r�}�뜄������"�ޅ鑻5�¡����fQ*�;�$6���`k�X_��/���L[|�����آ��!��4g��Y�/�����1�����c��A����h=,ݩȸP����o3M��۝Pة��M�.<�_�=��\6)��Zl^��ҳn� 0.� ��o�jM�����vn�s?ɰ)�d=a����$�LM5"�"��r݋�V#p3i�o�v�̥�pf�%�����}ot��\�r��h&"���Т^C^�⿍�Oks
[�����E*�~�g1 ǆ))�l�-
��u
��R��ӬT�&����2�s}� @�vC�4�sA*mFȪ�i�<����/��F�*a�j"��1^�����_��m&��
ъNm#��1/�kfF̑�b�[{�����i�؋Ԧ��Wy���Ck*�Y�<}�m���E[���\��POB�0W� �w{M�Б�T�Z��
۔-������ߊ�Z絧2�D�;���Z����K^ģ�H�=�B󇅺b]̀:�a� q�:��b�ap?۾��r3���'�%��[D�g�"d���9f��	ըV
��a%-�m��=���jt�#��\G�������y�&'O~����܂|j����{h���w�1v��Æy.��8+{{$"?#���-ڍ���qM=`��2�(�睹Q�rXF��N��v��FW���s�՟�('��	,��1��M0:�<���]�<�)�\�*�h�~��&���&�M�)��3��I���-Sݭ,,�����Sm�_�����i̩�xtn0��7�+�����
�ڱ�����l[� �0(��;=Q1��l�ϴ�i��X�7��������'�&�D�y'E�wl����3�i�I�=�jF���E��ms�G��E��V|�ɠ�����N0��w�Uk�E�� ��`��.�m~v�̚����V #���q�8]����&�����KYJ�u�<����ŊG=��q��bPKʱ��t3�q�x�����+��`��} ��+웘�X�ظ�����HW�m�����\�u6�_�2�Sy}�#�d�m�*�ٶN����{��^^ٕ��)�a�%5B�kH)��M�s�]WE�NFrD��\;�/1�/��"$�xR=�m�ȶa�R���r�g�E���h�v5���\�:_ϛ4wѫ����<#W��}j!�tlD�՘G��8��~�S��O�����Y�̍y)Uwh1|eE3I��'��"4�q0����S��%��1���ܐ��
��bK�V�䱃�X�8H��%�jE���j��H>Gkʬ� ~�Z��������g�������xK�$�\�oچN���vM9�&�CЛȄ
��������6Io��65,�܎U;ʍJ�^֢A�m�f|��7(Z�goO��9�@�oΖ�- W��'�l����;_*m N!$4��p�]���n��M���ؑ�m�wi&�T᫢P���t��!r�
]/�5��TW�����w�D���F��q��k���0�V��ѭ� {	n<��\+���6��u�����A�3;3<.NCt�m ��D�9��A/�(��N� Udj.�иF5Ao-�H+aj�|�qSТD6 �Zi�m��-��6'�E���V���K�v3j�ߢ۞)��lб��I����l�9@.U�8����8Ɔ׼]�*�k`��F�85��QW�d�:�Q����uCj_��5@)�?�^�~��8twN�o�:����)�P�]l��"�
��%m�	��J>̿L@�<۾����,d��Pm���,����"�0�-�����l�5v<���B�抹�S����9��U��d)�nD��Gr�k���"�Ă�1�$�mp�fZxo�WE�@�Y?}�G׭����;����TYX+���uw_Z�� &go��
>�K%���{6-�韻ze$��4''Q�̙/�2Mw�T<�w���@'SH��Cyz���x9�@_v �� �$&�>e�Ơ<=N�>��1O��H1�����**�z�{I�&���\�θk�9'>D���dm���wJ����=4�f:�=�;��7*�[H��4����I~L&"�W?���<P�g������y8#
 ����q3�����:Y1zc:-�<����<�\�5' AX,�
�dc�A�@ϣ�X5��Rm�ejJ�m:z�6�Py�M%��e��7Tj�^H��=�Fg������(6� ��S���F������x*�Pc��Z@Y��l����~ء�+��y�?�C���6�V�aBtS)A%�rWG;q6�P8MKp76E:�rH�������pĆC�%�^�J����u/��Ӯ)<��D�v����뎣�%��R�3QI�V�6��ȥ��Uq�&0C�v�����#=���h��}so&lt���_��Tp���%��e�����쏚]�Y�����V�㽎"�0%#�eB��A�G����U֖�BM����@��V�,�Vl?�kEV�	-��I�]F2��-� U_Y���=�BN�uA��;��`���fg�ņU=ű-<c4������[���T9I�wE��4��z����O�B��Z�i˗�e����'��i�Y��)�tϲ{���`ჱ�������G�R���0����`;}�����4��=E�݀����;���*6�PS�(�R��Z�	�b�e�q���xg��C�<{�����Y��k�n��S��j��š1�Hh����1i�|���(�쁟m]�#�)��a���;���yO�0��'_����	U��o��Cv����浪�H<o�(\N�@��0)��)�l���b�
J�M=��-����X���N_��!���K}�����T��镾�xAJ�YQ�|e0mo�]i���y�/�xT{,!v�*j�4���Z���� ��]#�� �-��7M���ϔ�L���^�� ��{�i@�!����'��T�㢪�ր�6�GxH��!]�tbϗa��S�_(��Q7h���*m��w)��q��eӿr��A���v�����03�6��Bt˦#�A��Y���a�+� �<!�h��nF5����Es�k�I(�l��M�q��l��i�QI/eNti}Q]6[���gb�^�U�ķ+���Z�u!�6�wm�c6/�q=�^S�-�^߹4!UA�c*��O�=~���"u����:���q�������e�I�(�Z��A/Ž���A�c��:������Q"���M(5g�8����M}��+zؽ.�8�e�*��K��B.��kMJ�
>X�F2Z�br�T�\�w���g��_���K�p�R֌>�y�9��c�����h���7&�AR��=�P�z�o74���m�{L=�AWq�L���;�6F_ � 8 ����t��X(��IĄx�maۿRd�Y|Bݯ�:��!�T��-L.P�d�R��tӀ(�.�ț�-�I#|�O�"+>;�$ev�>� wC[6jw,�sk�__|y�pȩ�Y(6v��\����@�ĩ�c��'^w��Y���KT�:
I�Fm@RO�cd)M����a�f��(ë{x��z���h˃������s�:7�m�[�-	�v�U�i��暻S�h���fC33j��nGo%"3wTi�~�ѲZ�J�og�5��^ȶکJ��s���c����ք�,x��{;���V�����α��=|�r�f�'�w��0�+�sl�fpY�O^ʹj���:�z)�����y��DI���c�L�Q�7U=xxY7�ڋ ��h�9��\��\:�s���N��N����n/��(B��/=Ksx�;�Db$�R�,CO0��S��h�
��y6P�����c���@���g����^�5����,���Z�U�(��q�x���@B@����0�&�Gg��_#�m�,^��-.�G�/}#��%<�d%��ք���gg��k�AKzk��n�C�I��(x�<t��JC��̜z[��^�oǈ:Rp��)l��͉��2'���gF�����׿�D�d���� .G �z���濟�̎�{[9���d
G<Nc��vv���Q�
�֞�N맒�:�Uh���c���=��ӻ��$�Eً�|���D
��A������tށ�8��E���Z67���Պ`"��}T%3���͘V#TǸ�u���n�3�z1����*�]"�O�ՙ}�X;�w��k�$�~wx�>VH'}���l5����-TP���ǃ��2����@_�4 ��^�JI����pS�K��:4F(����rd�E6�(��G���7]�fv�힏eU�vd�r�1��e_�$:F�R����]��X������[s~��d����ky-���P��3��&�J�N���[�uDAS�$j]4��^ g���|��ד7�L�VO���f��y������r��j��
���9Q<X&D�Kuh+�5�����x�P�̕؛�RmNsa��,{��������k��Ep�/wJ�<��cmy�D�$��?�O#�c0�J�1���#k��
"j:
.>���'�̈6��F�7!�yG7,A�@��V5*M�j�$�^
l2�&<[���0�,h,�O�RPY��n�`%Y�W��#ƞ_�{jM��%}��y���ˣ߹��U�ԲQ�[k�Bow�ڻ�9U�w�,-
��c2��?��s�>��IhQ�q-4=f���j����{hkV1s���A�ۊ�e_��?�rm�~XN$h�hW@��X���'/�JM�8��y��KK�TE�!�G�2ע+|S��ױ��wr爘�X�'�V=x�5"�lOY���o�������a��� 
+�9Q*tW=��%Ĭ��b�.I�e�+;�Q'�9���t�wrZ��-vH(��a_�i��҈i�9"1�Ə���]��O	�"��܁��h~i����v�{�k�j�G�D2����ݫ��xλ���1��K }:n��R=h�.�A������"�U4Z���a��>0�׺ և�Pd?o�W���%	At.M}���.�u�fs�G�CG���10^�-��lԨN�K����;�=:3���V�X��*�|�eq.���eki�$ ́|��f����|%�Q�ݍ�_>��j�����:L�J2���L�(c���M�?WΞQT0�f�y*� ��?n�P��W}Y2�|ホ� "� e;+k���H�gT;B�Q���^�r<,�V;�Ԍ������sh� K� u&��	J���c�o���"��Z��Y�g��4��l��F^�U�s����8G>i%����D�LP��K�ƎM��s�l�����ۏ��J75����N�˚v�m�O�Om���e��y��_����1�D�[� �v�|ZB%;� ]e�ͻ�i��נ^�隯;��,����˕4�Cn%1����3�`W<׎@l�SU
,�b�k84,���z��%�gRi�s6h	l��p�m�&61�Y�z�4�n��˞>����U������kJ�Ʃ^�����y�x�h,�l����B��6��b������)���	~�z�t�|O��ꁑ4��r!�w9w��+xVɋ���F�L?)<,+��!j�Vm���ap�)����ݧ�t_��n6{W���_	4�D���7�ޝ]�g8�{�gvqWa"A�u���p�P.�c�V�a=�q���X��H7��k�=��etR��/(L�b[-s�E��W7�iZ��,F:b�y�<�W�'>W6zj��iE���i��[����{0D�l*�!��H�78����4"��3қ_��Փ+�ٸ����U��u#Z��6~�#W��0�%WJ9��H~#��:��_M�	$%Ƅ˿��ʣ���m*����,t��t�1�"6��uY�ڡ;���U�=�ds����f��̫-�;�!I�����Ka�E=f��g
��	Q�`%D}����y�
̼���`Z�R���ԩ���]��1��I�	���ں���iڃ+u$�o#T*�lH��Q,���p�{�eR�^���?�����7�j�c�VL�a?�[�k��s�6�c�J���@�̶���=�FQm)�_�Up�����h1Vh�(��ټCr�#{�nMki��{���Ţ���$E�wE���n�������J�Jg�EO�����у΍"��Ӆ<�w[vZ��h�w��i�1�{�o:�T��;�R����:Ja�0�l�`2'���	��6f��֤� ���i�9��|$��p\MmEY"6��3a�p�7X�ơ�3��%C�RZ�M�!��俚��nX��.�P�U�����\d2�D~/�v!l$ٯ��V
�v�~ҩ������	6�9��a�g����}���"D���)}�S�M�r�'e����}|4����R.
���*�����*�#����Ϻp�8;1���p;�W�<���>et�*i��h"�a�g�s����/֪���1Iv����$���-����WȒ�>-oi�p�q�yuX1���:��&�l3��Mv$G�	��})��k��QN s�n�����\#��-L�W��p�IZ����X�G�؏���˞/�W�+�-d$�/���y;b�I�س��	qک'<U�����&������:��HU~:,҂%/fG��ڠ�E#�n����觟���QA��ٔ��8
��\6�(�M�Dԑ�1aDex�׽Qxn�GȦ��d%��	[��q�������ŵD�� ����3���L#��7��U�+�}�D?9��������|P����&,^nko�g~����a|�g���4t��.�%�a�"{� rɁ��ņ6�د�<\�Q��Z>�B�q�#��lW�b���"�{RP3u��%/ۼ�$���Z�v��YOkb)�1DxԦ�h���26{~�H40WG����m8����hl~R~�xav�^�~�K�`��H;p�]��i�c��m���3ސ�K��i1�����9�w�ߔU\�'-���z���=)��D�/�Iqr�ְ���-E_u�\YMN<�W�M�U�[��g�2����r:�Òs�z��H5�+d�:�ά��uw��@nÆ��=Ϟ*��+��7j�!<x�E�e~�Z��=����0���W3��[O�	���?���Z�D��!x����`����$`�4�oi��:�$ڑ�y�f��@p1����LRF:1++X�`�	�����@]���u���^�ϡ����[�+���8����:u�qL8�˅������s~��Z�lOgD��m_x���x�1�V���P�����Us▮x��Y�����Ĥ~��X�p�N{�5o�.M��bm�NU�ؽo�Yx�X��U��7[���%N�X> p�p ��b +�s���'��Hh�;�70MZ]E7�Z��^kn������-:~⬎l;l�7�Z���z$\t3lr�ZD��fT�mu�#�t��;ӻ4�����^D_�s�{)`��� �Z*H��'�RBk˩r����'>J�0�t��M��SܚtGԱ�N�,Ged)WCN�~|+��j��q!�S�-ְ�}غ	�K���\�W���.CKZ�	��g���Y���W$X�`����H�)��\��_��T�g���j�H�`�w�kX����L���?�HS����k\�uz����3A�D���A;zM�DHm�r?|nKD��7_}A$\���)=�9�`;w��n�`��D��x�� �
D)2B`B�y_L��v����h;��-�U�x�ܔ�OS�cY�^E{.��d�F�&��7�C�+���Қґ��m��*�#��6���W�!.��4�lwN�m�a��0~����[&����V/��OB��Rٔ�[��l�}D$d�������dq3*�.wk"RS����)Oys��(���&�J<�B:CV@�
�������2�(�+k�Q{ۑ�0#��5D��lӢq�o�]�,g�!/Z"c�[z7}���4O�B��q�k�פB4ȅ�UⒿ"P��i�kT8�}յ�j-G���<q��M;��	Z@�IF-���w��.��Z��P��~�%G��jH�q�2�G�"��5�^���]�l=��sW(^�!����pnm�v���hˑ��_S���>��[V�m
ȴ_b�&
�m��l�[�x]�/��~�҆�فG���.��Gq�	k�%] ]TA����TkE���2��^<�.H�J��U3���+,�FNU4�"�>��"�%���3!�6Y9��kʫ-���̱���Oڹ���ԓ��W�_��rU����0J���ڇ ��q٩�]J Q��= 0"���i�lNg���*�uOn�`J�"=��z��o���K��@����*�Y��)���G�vas�ӽaZ®��(΅�_�2 ��������0 �GTc�ޘ;�����Fԓ}��o<,����7�>�H;BDpܣ�W�O��<��)��'�s"������\wW�_CR���F�=�\���PZ�}���>?�;P���2{�U\�d�k�A����I��Cz��ʱ�VV�Ӑ�Ä�?Q< �V���&n.O0�����ݹ ����B=^�����U�E����sS�8�h@�O\��:_��5cf@O��nj����������t�ތ��?F�q8f2��J v�_bՇ<,}F���F��
P{q��9�]� [��t�$��Eyn�LmKAF��J5���<�us@\�F��=���3M�*��G��,�S���-����j�����Dl�l]�?Ɇ,��;z����I�BJ��~�X�����T
6d��Lv�E�i�C����2e8�=��։[�.�~�n7�O�'O�&FN`�D��1�Z'e�N��c��ɛR/��p�b��x?/� w"�x��4�${`�:U?�e�W���6��˽�1v��Y��'*n-� !��F���Ʈ�u{��S�-AXeu�ʖ�������y&w�Շ��STV�����NjŮR��s��8JmvE����x<�`�2��T�2�D�Q`�SnC�}����eY�#�L;�=�[}�I��xM͘��~���~!�~���7��X�j6.�Dj}�TYҰ�<�d���h@X��#R�Y���!m�(�y�ص�?[b���]�`ir����$�^�� %���&�t�n,c�L8;�u�f���s&���'�Ң֮�.J��Hq(��T��DNTf�\K8I���FL�9��s_���`�#]R=X�V�Xġ>䔏�yf
H<�QE:�!9��_�'B���3͆@a�z�8�D��9@=�U��Y{�P �׿����f���p��"$. 	l>��1q��G����u|���]v��Z¨��S̲�=��}�gl�[m{K1�1߈I�p��ʛeJ�x�=�jB�*f�h�!z+���d(�H��Y�H>���o"T�- ��W������t/�#<$4>BZ{k4�wK�'ti=H�p�W�%1�h�����fH&gڄY�����!�ri���!E�;5�QwS�t>��x�(�ze���B�e4�cfJy��Y��UI7�R��
V��ml�>O"�S���Q.8�a.U�Z��RO�	�}�}8�h�%-��Vw"��e���7cϼ@�F�;�m��.ǿb�Z8�|�0<��G\�^n�˯r� N���K)�l��AM?�]��� p�e�Jb'M�s�p�:\�)C�1��p�4+��N�q#��;g����qz�6��(�h{ o��j��X�@�� ��(��5K�}<��������}�M��0�+ [x�RNy�����+������a	�(�
>���s�_���8�����P�U._�Q�����}A�b�ⴳ�H�u��U,bX6�f��l�����p�d�:�����y�vͻ�oT��K7�M�밮�AtI0������?��>�B�k��(Y�X:�)1􈏃�H$!+aS����rⳮ�@(�Wm=�ԻL20���Z?���{S���V�F�_�^+���Ʃ ĵL��3�5�P�Y�*ۛ΀%��a��dvv�.����T:z��`�_�K��vl�|��� 덽za�-�J�CC��,�| ���ϲM�Ta}M�d��6��jN�}��$z۽���6�� +2����1�t��e߾������-*D&`W�bu���Z#��Ɏ�3��}\��%x�\	h
e��ͱ��D������y~I�&L�2���P���.~*%]g�zx�m[Qg�$����FkX|C�T*̙s���H�R��sI�l�b5Y�����,�W.��
�N�v�mlj���L����������&���sD!�C0�S�TA>r�|�$��{m�ږ�����$&���61����2�����	p&�uC`��l��@�LB�����7.���O[?um�VR�0S�7b�n����a�R"�U��X����&�(%��=,/���+�x�f�;��n`�[s�@$���Y��ہm�c�\,�b�C0�J\ھ����C<����� ��!~���V}ߋ�Ԥ��3T����1�J3�Y���L���,�x�8���h�Zֆ$��g�6�.��&�����W�4�Z�y�D9�[/D@ ���9�i쏡bvOD,ڍ�!hw��&�y{Ā�}c!\?���G�.Qv;�ɿu�ܾ
�#�k��X��(	�jl$j,�P�tzcؽR����0&�j���Kc"U_*(;d�(���S����cG�Ծ����iG�����V���M��Z��5��s(:{��m�s>�-���/��~׷�{(�?�����4m�̻���?�r��Ӑ�T����c�|>��0����xgx����M�U܀���s�;���S�����Ƀ:f8'��Ƶ��vjD�4�D7!@�X���X�����G�Sd`Mk��

���/7�H�ӡӸ.Eç�rb�P/˿"t �E۠�8�a�!/�}x��s��f���[m!��K��0ћ~�"�O�|���gW/{_nVk$$�.�P�R��5sZ����v�4�/�}��
�UF�{�`;�Q�ku��v��_۷诓Y\�Vd�����W�(�H랪a0P���4�u�?[V|d�x�m#s���Ӫ����D��<�_��!H�bTd8j0p�ˊ8?��Z_U!���X�"֒y�iM�Jc�ӣ0�����\��+��FO�W잍�����,҉`���i0Y�C�����D��n�<�3g���((�de"Kw����_g�a܁^N��]���4Q���To��X��#��q֠��*�X�}�^F�y����"�x*:!�ycc�oH����"m�5�
[M� `�Q��ƕ�DS��̕�c�M8��%J��*������+[�񔢜S]�200L	H����my�N؃�X�m�f��^L��5�G퟈�7�Jc��~
��I]uy���ߛ�^��C����E�dcگ��$.�H�ɕXF��.�|x�N�2NH:��
��m__ 
M/�Lr�Q��c��I�I2F��dR��|��"�ͧ��5
��%�c���1y�m���)��˴x�K�Yu�Z�!�r,/���c�P�;h �Y�.EGO |h�4�[tj$���ub��sc���;���B�4&κ�P�ۗ�s����a�uy5�a�w]��o��X<�xꉟ��"WC������/J�cb�7\ �_Y<x�t�X^Eo`��ȳ:��d�
�Vt�Q#��֜�C�	Q�$�}��ҧ['�A!��Iʘ�M�_e$s������5�+J�HԄ�fO��
	ɰ:��Vb�l��)/J7�u���IQ+x�V]wI8���\DGΡ�Fn] ���.��[Z�Xlcs�Y����� \Nn'��̰��~� ��Ҩ�MP�*Ѡ1������0�����5R4owTR1����h���[�JHom����@!qGI�ߣZt[qU�w�i �[Ö�s� q˺�MCm,��j����o+����`�up�8+��l��i���՘)S��f�����m[�}����,ňm�mɻ��O�T���
��p��� "'5�5+���'�hӔ�8DK*!/������K���Ѕ������i6��]u�,?!������\W�����?b���#6�EQ�XH���`�����ù8F��
I��$�XY������wp���QG#J��o�CO�N��/�C��⏓�.�������$��߷������g}���J�����m�M���W(�������S �
"�6����Y��q�8�H-�I#HL�K|(ö�v�v�.���h.�u4GwG�L�p8������ؒt��ޱ�F9��z��H�A��y�a*x�πu�>�@�oU$���"�Wk*k�w����nN����#z����Htes�Ѓ1|:�)��e�%�f#ź�%���)�P+<t�� 0�E��֧o�ɷ �#�"Y�����x��:؎!|D�1O��s���r,Q����
S
�HZ	�<; ���k��!��[;��j���_�T�*}ҝ�m4����H��׏�e]�]�8+
����P�v�le��鶊ۏ����m�D~�N-I����ޣ��ν�f��X�P�[�#m�Lm�^f�b�˾JF�y_�ar�n�al����z��a���	��	�����"!�p糉��V\h)��*t�MI��x�5�KJ!�e�2ZO�B�z&$Ŵ���?�����Gs�k����V.��u�a�}�sJ�nu�n�QT���� ����֢F;���>�<	�TB����E�֞�S@;�pvݣ�x� �L_
�z�[~gv7���4���
��(JZ��3ܑ!j�K�� `Cc9��c3y��'�)ʉ�\����p~ozVq��Ay|�uB�n#�rL�t��A��$THR&&p����p���%��u���̄�� �5\h��@q��P�N��+ Y����'t]>�&\2܇f��y��A������=:��_������O*b�3qB^?�p��xe��m<'R5&��0�:R�CӁ���)}[�X{nu���2k�}-� ���v��Ur�z����kl�0�`i�@�����	��|�˿՘����-��e ڮ7��py� �%= ��F��1��c���1����C��, ������ٍ���B���e֥,<���]�����G�l��K��]�F���Ja@����YW��C�^g��k��v+�u�?�KQyYMc^,T�"�̾^ֱ�&2���&v��O���F�q��� Seu2	�����؝n��T�4�L��,�])+��A���r~:�@�_�f*�Y�SW5؊W܂�w�����u�EGG���O�f>�dlS���^��W$d��+��V2h���y��C@\'`ԗP��z�$��M��s�A�y�ap+��	7����"k��L7t?�˟�wr�xT��*nBr,��J���6�|��9�[#�\��@B��p� %A��H����ی(��5����[�F�9n���vA�5���Z��*�џ�kq�W1V,'.�T�@
�7;���ϵ/(��U�]t�ݵ>D9'j��	g�ω���ۣ�ek��~p/�+�F?&��л���﷠b+o�O���%����=?��ZN=e�#L�-�Y3����E^�zt|h�ï��E� ������6fɶc����!���@����l��� rC�����ֱE�����8��i�,A)w���_�N)�V�ȶi���y�RUQS�,V�VI��=:P*9�E����6�'���0�|�h��a澽�tP>���j�Nh�|��w'�ҡ���f�%�����ZȖU������������"v݃�%'S�5t���X�:��ՑRƬ�ū���J3Hya�eDm�
^�/~�{R�ZP*�	�\�G���ˎ�g<
.,��(���bK@�
ָ8����"{נk�D�T?��Կt�bsl/��_F����z{��FwBH�8��"D�&��q7��a$?v|a���,�BTC�70�ZE�<X�:-嘈��3IP7��Ur� �8��AvS��	���i��wb�^����+H�"����84ܳ�r��ת[�z^%��(W����qa݉�d�8�l�����6������0줢]ӺH�T�����trO�����U�w0�d ڿ�\����:U���]�U��䜻W��[��Y����L��s��$�;wCV%�ԙ�)D��Ӥ�:�ƼКc�)�aA�;���]�if��S��;Zl��6��V�_z��}Z��E!	
pN���G���v��CĄn��]�g \�������q���5���a���Ў֡;pC/�"M�c�o�F����9xd��6���Ύ���P0s�Z.Wp���9�_V�O�F\����~9[����&������ؠ�����@�w���0,{�`��nCo�yR��`Ad9]D���H�N��Ìe�=S3s�9��C�!�<����r���eFR+@3���	>�F�W	zw�[b$���iE�I#o��1�ߘ1F��UFn��{p���V�Pѹ�*.�)�?��%�6##:X��P�Q�5�B�1�'��X4���qp���xY������+d̻�b��lL�k�D��c�8'�����Ȣ�:�C4ի�Ɣv}����m3�T�t�~1QrF@L�ެ �M� +91�M��As�[O+R��yX�7� �� �*��P�$mgxap-S�ay�����xڪU�0����A���0(��P��I�0�o���#��dL+��+*������F����|fC��j���|��kf�]��`�L�C�@��o�o��함v�U�e ���5�����V[�~[bbT��<��=/�G�Xu�g[�M�������P���]�`��oOl�i�f��������K8o�K�0����kĝ���ɷ��}o=R��K���)��
��P.� P�-K�z�>��Y�\���!b7��L�f�ڟ߭�PI<�R���B�z�h$`CqU4�Fu.������
/x_���Կ��*�'���s� }(Ԥ�Z'���:��N@�(Lji�6	l+��l��M��M��w�h�d���F�n�u��,Gf[)=�/���f_��r����d׉w/����5k�E�\�Y����r�:�LJ3�:�ΎPoհ�"PyF⸡z���&$C��pP.�����M�B�߿uZrE�8�m���<@uΌ'{�����,$k�,���Ӵ3Y�BZh�Z�;sFx_�Ĺ;�P!�L��z��xZO[�
����A�BѦ�)��EO�˴�Ʒfҳ��̔B	aǿ@��1��0Vi��~.��߀�x�l�A~���?Gq;ú�)~�2
�.������U�L�l����)�e���t�'BqV�zK�ՠ�/7�ڊ}���;^��ǳu�O�>ja=�k����GO�SZJ��RX��d�+�z�	Ҡ\���\F��zn��K� ���8��90{�dwR�(���k}c�޽�t-4�@Ő�ж�0�l��i?kj��nl�S���ݒ�e^����ZǵM��l��(��jh�ض����g2�_�N����Au�5�$|��ja]񥍥׈S�e�?[��Z�%u��]�c��I ���tM-0��Oܿ����P �a|3��s�sR�t��ow�tnƷ;��_��B��{GО��K�b�p��M{o�,M�:Ib�7����ƨ�]��g}\��E�P��J�q�$�,jb���N;F2��V"� �ׯ�&c2�e<u�5�fw7OV�MJ�O��o��������5�Lݘ�z�ᜇ�k2A � �d��q�:��0�%.#]j����͝,�/_ٌ�R13p���\�k+�r�BWa��[�*n`�Ebk#A<��;��#�*�GK邍�VP�5��ƒ$���kU"$o�4�b	�UWC�!$[`��w�jL���~B��X�U�����";k�"[Q u>o�����Z�xnB]�E�\,MɄ�r��Y�g��jH%���n9�k��}V�Q9�w;��-f�W�KƦRڢ���H�� �; j��̿�$��@'@�ԉ���S������}5�pT� �g7r{a��
�A���= �)��7��Iw�`�zD��,�ãg�� ��� j�����ȔRv�`i��+Y���v��93j��B�������$K�y��6,+I^��6=�t6_]���iq�z�) D���3���?�k��g`Kj' g���J:�Ce��D���,�Ӊݫ��>:	э��9�@���[�䡌�#s����r���PL��7��C�?�����H�t�}��`�P����H�{��`��=Y�)]�0��(Mt����3�і��7�l%%����c��s� �����x+���S�L��򿃐���N%�.����II���x�����5qF�e�xP����D�������5�Q����DZ�}�Ԁ<;�7D	U��jq⢒�^ѬG���S��%�;4a�v�$wn>6�.H�♋0Kr�*ԓڢ>����m�uxtZ^��j� �[dr�����s�kt3t�PK�K0`Di��}V���A��q��s�����}.Bϗ�16p���S	w,�d6P�t��?�\��]1� ��P��ǘ.o讴m6M��X��H7_ۃt5���9�ёnf&���FK��Oao%�8�m�,;c������� ����(HS\k��ì��vX�8)Ϡ}���-�W�A�F��j�2PrX�"�.��N�r�7��˔�d�p�ӫo��޶.�r������A��9!��Xh2�����,I��2��P�&�I�Ѕ�&��M��K}�<w�#���6P�[���*�c_�J\'�k��.�3���}Ԗ�y��lR��Co����ws��������@���KPAh�ͽ�F1��/����Q���#��N	��o����FK�� JR]�`I
V'��[�<�+e5 ���F�k��8�r9��-^%ñ|Y��xe�#�y�Ys�����A��%#y ouB���6v�v��ۂ��7��&_pmSDt�bݜ\����<�s銯s��fG��X̾����pESr�p[����pV��d$��,�0�����-��	/��M��\SP#W�}���𺇷�/`����fN*y�+4����dx(rn(��V��_3�h_�b������Q� h?C=���
xٟ����r�f}G"{�R:(�ub���߲3�:JK���<��ǥ��;I����_Z�	kbD���)Q��y|z�#�I?h�~���Vt$��ܟ���Ɠ�ނ���z�\�i>��&Ƅh�N�]�~�-<�Px�rĨ81���������C8��Sͣ�2�>�IeJ�j�"פ[{�2�3��c�ہ��)�,<Ʊ
T����"1t�Y��ZsT��8	�$=�n��r���
}��[���W�2�۷h&Y�_L:��>z��rV��af�!����V�G�-��@Pu�@�ז_6�w1$X������3,}D�����RJ��N���xR�^�2�ⴛ:Z$rW�
8�ߟ�Fj�����V`9���dn�	�t�Z��N�`��V۱Y
5��!f��ܞq�@F��+�1Y�P����!��ъ`q��G�k�2G��pMM����zXo��G`�oB.ͮ���`����̞P-�2�s]'nivN[�k���%�2k���Y��$�7pϤ�-��n�1'Hg_N�R�x C��;j��\@��c@4�87��}�y����o�����X����Qvɻ�ѽ�cS��6�y����
�����v%� g�g��C�\��3��;+��#���[sLS@��(�$���K�� K|�a` �c�~eiX��x��%�>���D��_�K�pN�[o����x����$��T[�ZDy�Q��L_�3͐=�9BaЂ+��]�ȍ���Z"W���+�� �Hx�����N��]��c��4������^��}��Q?4}����`� 6o��j|@\�(*��:�����Z_�.N�>�)�ut���hmsu�!��k@?Z�~u�=C��������z�<L���		�*���E�"��+{#��U�5�
%��.�g�4���6+�rYj�U}��vMB)0��ԃ;�����b�p{dW�k���6j�m��o�����K{h�t��xg��	j��H��s-R-A^s�� �����V5/��6ŏ�<��I ���Yh�7��x�J/��C�w�C/ ��J�
=�9� ���8)���m>R�����ְ^&"C8"�Zb碣2rI�y�9<����:��3k箤�TQ�H�!��7��l�H^�������Nn4Fޞ��uFfX�[�*���1T%�6��L�^T�գ���xԻ8�噦�w��n���u}>q+w�L2Spyq�.Y�U�{g��wi2�/��
������&���X�J��V?r�j�����E��`��c��`�tOé-�R�%FT�a�T�8l�{(���@�t��F�~E~��?$p�zCG<a^ ���4c�l)�)� �C�wd6R�\F����O@�����7'�Y�<��Tw�^Ѿ�||���_!,;������ZC�s�m�>�~eu+�h�I^�����DH�f�c8�4�^DJ�֔����)�Q@��t��Zˈ.k��O>��i��d{Y��{��1�2�Rc ���%����]y'��]�n�^�<�J 	������_�s,��@�*^�E������T����.���	�������a��,,`�섙t7b�0�⸈H�ߠ��*�����S2��y&F��U4J"v!U2�`|A�X�~�����0�*���?9�ӥ���s����Ј���(�u}����R��=�ăH�M��T�ϱo�Ee��o(��)b�a����:�� #>F`v��m�D����5��Ӫ���zsN�./O����UQcK����խ�C+P�"8��E�X�4��bf"�JP/<��:,���3��j �\G�`��S��0���t���]�jKH��)�t���|�`Z��FO�-"��E�4���S"M����(�S��H3�.�I^�gxؾN.����i=����"����dRV/͡Ho�,��Y_p<���i���RScI�a�'�{�61��k�eP�'%���%�얀s���B�p~�$����*g^R(Z��	�}]�.	si@�q`���p:w��f�d�D5͕;��H�xz	�䃐���%�i:$��(��;M
\�����Ճ_48������1�;,	�I� [�������YX8�̿�=3���eQ�z=�:��D5.��r��n��U4s�u��M��PK��Z�:�v��Qѧ?�8�����{0��:�x�ɦIOɷ���r����h\(*��	�~dM'��Bf�L������� *��Z0�FRS�fPzW��Z�6�"}b����2TG����j�y7X!�=А��{��FB˕�ɚ{4�x�A�G�~��DxP8��ˇ�8�W��I���&��#E�(9����#k��q�|MB� [�����ݤv
S�9�̄<�Ģ*a���'�"�����v4�ID*��O��!�t�UW��Y��^���ݿ���F��H���i%�Oj���&+SL$-ѻ뙩���jP�����N	�E�T"ĕ1]����ճ��	u�D��iad΁x��x��B�aL�a)���%cHȥ����d�<�$����P�a��_����u��f�a�l�8`��¸�L	?���uqȤ Ie�|��4��⳥oM\2��w\����0�)Ğ���Uס>��j���@٨t�N9��Q\L�>P�[Ȭ3�pnT�r����n��t5��ԛ�ھI���ê����3�����:�yT�v�c$��~;��A��32��7�u��F
͓�ls�9�y:�8q�{��JO���za�������(�^�<%h�(ẽ�0�2E�ܓ�O�{�;�I���<����X��b&CD��QL"e����&_�,3���	s+�kX.�r�k��?|'�կ���9� 6�l>�`G`�؜�����ӽ��.��Er ��b��A�hܝ��J�ˆ�e�Yh2w��NQ�&F'��Wb$W��˱�|\QG��L.����tZ���u���tIw~�*aT.$��q���T�P6'���JI)�a����au*wo��\�mU�K��D�nV�N�A����n�v���&.6b	��z&A�&�Q5��o�܂��|�����N����#��ʮ��Ţ[�`W-=�����O�2 R�f�Ѱ�h�Nh��m�&�,3.<�:���0�Zk�¤���.ҖU�8_Ku/{:������W3���no��2��W�ĵ�����y��CynU#�(���
����W�}��IY�!֫�{�MD��X��!E��;=8g?��_ό��Cؼ+�s�I�F1gB/����$�����$#q��i��hV%�Њ��L�����[��mIQ;��ి6;���@7X���kOaS��:1���ͺ+퇃����Z�g�����QOw�?_5*\��S&;���0+Ń�g'�>o�b���{8����ۈB��B�@n�8M�4��b�fH;�X����T� ��u�PM��H��o!
��*�]��`��G���̡�*��	�7�v�B%�����&�w�Kq� D�m]Ƃ�V��$W[q|.�g����A� 텰���Q��1�-�,ۨƦkE(K�u0e�H�+#7+��C��>&��Ws��.	��ޟŧ�Ps��apg���)v������na�3%��7���z�_2�Ў-4J�ymt�h����pD��EU�?�:���tpu� �I9#F��L~Jݪ�Pmn܄�w�O þel��Y���
�{��X{$�]����z����Le��9K���H�����\�M�{�򶦫�D�VX|4Mmޒ/�:"}͹�g������ R�.�*�:WIH��}O��z�����H�����Üv�e��@ܨ+b�o�G�ͭ�Fuf������(�)OY���C�g (�C�[L���7��F�{*·��΃�y ��l�W�N����h
�V�F1lL.ox*���}��:ȫ��
��h���ʎ��#	�}�%,��P��N�a*t�)�$9`���)z�9n�b����"S�^ݿb(]F5`v�SPե��\~�󀕉^�gStڱ���%��
|�k��!���ŋ�&��'�KO�i����׭I���^|����Wתڨk��лLBG�6��K�-�`���x�
��*���;���K\P��j}x�},i�DI8��F�)���=Jq!�6�B���.��ZP��d�R�Q��>���a9����x���8��G��U�?'0��)Cn7�ⲣ|rR�����!����Z���%�m`���Z�Ӆ��,s#D�'�A��ƽ`�~��{HA0T��1��$Kҝ�e	5��-�1����������n�m�F��V��5�[�������1�>.Z�����ct�G�Cb�{�eM�̜'M�+�q�˫F"	#�j�ӛH ����>3�t}4�J��:��	�Khg�Z}I8.J��_��~%��+�3�<r��#�t-K(*,��z�z d
��i9���.�zRt�zNG�3��Wż:��e���َ��/ ��d�3|d=����E ���5Pz�=dq��)���X�\ �z�p^����Ԛ���| &��w}c7g�ՠ[��E�#���BҒ}6�m�T֮�����!|�_Z���}���������(j�^�בkӬ�l���.�R&Hb��g�����6���_jE��-�l�B���5~�.lU(c�H�Y�	�u���y�h����^�.^"x�d /�cO"�<[��>mPEӠ�JZ�`)��x<'8��f���轩,���1�kuz�]k�gz���n�4����4�T}"
JCM	9���<�bd���G2���v);����*i���r��P�s�;g6����P0 �7U��\5�������J����!OЪل6�]�MM�h������0j0j㍌������=�ַ��sCiI��xAb2���M΁�q
~W�xt�q���N���jV��(T�޻�q��0Ec��'A���}�c{��/X0�&m#�Ȃ\�3�6�<�3�����wU�_�5#�l��3�m�傧�P���e������&^X�Q���\�yd�})�8+R��5nc��/ᄹ�vx�<�`L�Y�����azI�U���k�{�Ҝ�%Ĺ_
�7��s]S�s�Nc���'-��~����k�M�����߸����m9Y^��눍]ZA ^�:�@Ď�M<Q�w���{.�e�%�y��G~��<`3R�@��$�!��G*�gߋ.^�}f�����mrNzV���,���in���iir9�����0��1_yo+��	`_ك6$x�게��@)N�Q
�J�-�Ҿ��EKP2��]�-,�%����� X�Ӎ�#R��h�;s���i�
�.m�3w��f0�	J���e�`�=�`7g�����2t�w��4�MԯI�enp�.X�	L_PT���Ր�PS;��~�x�Ğ(͝p�/n�>�����$oİ4���j8�u�o�Cǻ�3I�(����!�T{M2y�Ap��#@ۯJU�/�[/���c	YQq�i���N��w.���Q/b���0_w�쬖�!_��D�6Y �r��(����Ϲ�́.�ct��P}=G����%`�k����Y�.�N�:D2�r<��ϋ��t�>oٹ�QX�`qH�8V�f.O�����hFFh�ܒb')� �L.������|�!1���iџ��	z�O��"���5<O,����(�Po�xȣIv�ܺ��?C�h�HgH0mX��#�WAV�����z�?�O�܌����b�����#�?��ą��j�y��*{��EO}�5H�3�����>]�>�]qN�Gj@��s����S�� �̘���;���c���%W(�m7v�(���Ym�0!:bE�	��֗30�s�զ�8�'�ҠbXН��%�Q&lk�w��9I��Ϩ���lS������>���h<��;{@����TO�='� wĝ�r�B�^VT_3م����C���e�C+ %A�>��R������F��F�7��Jqp.�h��D��?Dخ���;���7����?�c�քH�����51���N4��p����-𔀗�!Iʫ�^�&�6�T�MW�9kzF�T�І\2�����l��&�>r[.�c��Nj��ً���S�͹?ߏfk_���5�w���/�Ef���N�ǁ�y[�y���.c6��t��O[�悧Jr�{=�}�ݱ�ڌ�/5��u,�����ޤ�My�%Z7���Ow,֮Y |jL�+MSYt=O�p���^c���m-��;8�vC7�o{�)��)�Ԁ�ЃKj� U�ߒ,��� t{�J���N�RJ.#2�b> ���� �$S�T���T����t�l��nm�,$��`]b?Pg$�w�j�:�	ԛ�JmX�\�	� 3����3|��Ȉi�-�zSf5�3��]	x���m��Q�t��j�{%}6��OP���vJ��FLZ�WhvG�>�9��K�Dg�m�$b=�_�+g�#,l-��u�U��rZ��i#���N���]��0��g�]u�v���q�<������ԩ�4�ߝ�n6�h0F���<\�|�m�i�����{���]�4�rѝ������3��Ŕ�W� ��NXzK�%� �`K�OV5��C��bl!��E�&Z*+p'��ϭ��mgk��Zp����-ks��{}�E��KL-�r���k"%Z��n�����K1��z��o`Wɛ�#�7����J����QW�5/�����K�j��V���u|S�$?잌0p�(C�*�)΂�U������~lK�0��Q,��1l���	�ε�s��Y~�2�0��Ӕ��/x��\�������/���Ɖ�r�g�\�Q��+a^3�f\�:_q&�&��_�+e�ǯ�cӺ�n�=�0���̵6�ϔ"�Jh�Z�6\�x�VcH��T� B��qĔ~���z��璘�"�/.��,��A��7)�t��9m2��wǋxi�'4����a3�ٲoX\'u�5��P�'�^��cK&��(�Էg�͟>�kz8������G��s�a�t�i����mm��^����M#"�g�i�6~ItA�F�*B
:��rU�QQ�kJ`x>~6���(9�x��"��6�ZW�©Ƽ��ǈb��l���5Y*Q�i(�w��1텖�qv	W����斨�{�K�vn�6���2�eA>�'��\�u����_�D3�`#��fW� ��M��\��v�����:Kf�1) �A?tM:1�}�E3hY}Q�0��+ts�#m9�>�@	~n��/�Ԫ�R����NY�B�@�52�B�+eA��p�T�%�1F�bb�d]}�D?m���@Sm��O"s��`z�H�,���f�uK�q:d�{R��7YD�`���mG�������Ů{�H�䯩 3�R�Q�p4�O�V&���gj+�4�0�9�|3
��(��T='Du'~a������:���6U���Z�.�p$�LS`������"� ����QTS�d���ޥ5!��`��ʓ�/K�!�r���ՠ���h���TE�ِ�Л�Gf��"�M.����[�9�g	���6���AF3-��U�+A�oѹm��>�2X��Xi,�w� �M�"��4T 'J��S�.���h͎3���RbǍ�M�&�A��.�n��So���G@I�*e�^䇞�a��ƕ`�@��ω7��O�>���H�5��S@�h�끡w<J�k��o�!�&n9�}���?�X��ժpύm���'��I�]:�4K(٪�=���A��3� �>Qن����f�ϡՓ7��)Q��N?���>#=Y�P;�g�('z�x�_�J(�u!����!���?p���C����!pV��I$.p+�&��<�!��{�[�\��� 2W�`�bb3�)�|��[���;��1V���k�|Bc���_����$���t6$
��Rh�D����$��rr����-�B���&O1�?�>�Q����#<���{ϒ�w*է��FxO�����t:e�0:sk)n�^���Hw"T����ʱU'�M@v!-f��^����ʬ������^����T ���t�����0�nȸA�����+��w�ݒr�����,MC�<�F��h�kj��͠4��(�1~DN�v9��s�
�ÏE��S:�j��j������=�D:BA�� e��F)���´>mӏ��]R��_��o�ժ��b����s�I	�<�t/���iT�S��5%�]��>£�����ɘ�e�`�'.�r�������hd����K���mp�N��)^
=ʁvf���|�Y�L �y9�	��z�\�Á��Z}S"��������x��ޠvK�2e���x�e� ��ԻxPJ.��Pu�U��:r����٣���Dq���;��у*Q.��0,�EI��+��Ot?zGU+��.I����A�*��y����"�=,9���n�)��3�rV����x����π��&���W<l-m�,
�����ߙ��v�/[@5��85�	fyB��F��{`\=�,�KE�⧆�q:��2�u�p�����F��qybL���#���%�<;x��>��j���O�Y�@U%; �>W���$V���d��$���5�������tF����(��Ns��&�8��ۏ��b����S���
Mx��DX�"�x�Z��!='�l� ��"�;Ψ3�OH��#%�PxF%>c���4c�!W�����:��mb\@���Y"chz\��g��a�s��Gxɣ�ϣ�i,�4(SM�ʇZ};S_�x���w'KE>'���>ݣ��Ʌ�+=]�R����Mv�4E"Θi(���Ͱ�ݏp
������)���u5I���l!�I��SU[#\��w���xh}r��%B/���]�����k"UBjĈ0ܱA]�	�/�9;1��UR������k��N'�F��I�rT��齽uC�Q��D5:Qdo�G��{N�>�I�2iJ?SҚ����+-8��tZQg�h0�a�#ߔ��� ���N��?�t����{�޹%B�'�w�0��\F�������A2�_�P���}ǣ�8Wg��ֹ�1�`*V��~�� ��y���N%_�U`����x�y�	�&�X����XVW��{C��		q'�X���p��Tő��$v=�zAz�Q�Q�1�E�n8��wJ�K�GK�.~�~w�^�?N;�5��9��=��� uf�o�Y�{��ک��&h��;��F�d�,o��W��fU�ItCtj-w��k�˹�?Y}�*计�g����%�p^����%�&Ccc�l�D��J���8&Ռ.�xE�d�we(�%�X`��!��t���8��������t��v@Y�ַ����^f�S���bX*���Q�K @(N������g:�WB�A�H�N�'�Kal6�Vys���k�o����XG^�in�!�O;�����R'��k��V��ξ0L�iѨ~�6k��*��M;��A$�d3^Y|� ��dj��cp��x^�� A!�wXn�5�����]�����Z�+����2y!	���樷�ԮD_ ��K��,�M��j�"�5#�-t���e��~C�@�q�=���[�L��A�fmԒ����SA��Z	���Q�"9��yp���<	�K��C�IeI��L��tj�~skRt�>e���y��w,���������E��	a$YU���(J�݀_����Q/��L��'&�|���,�$i-��X|4W�O�����Bq������g�~�C�g5��(eN����I����`�#UD�C�������{�`QA���JtKeIT��`!�L�I���)����
�g@�/Fl��cQ2�-,0�8��Ʈ0�g%�:�`@���f>?� 7Ĩj?����Q�e��6w4:�84�*Ҳ���}le=��4�P��~����A�A&c�q��^�xU@��sx�]1-�_^ҍ&�>���������Z��(���T�=��1��"��I}�+�u�㘴�0��%8E�k	��m���}�=ٽ:�������J�"L�9Ɉf��<��O����i�x���%@�R��8����Lc������y�S�=Z�Ou��bS�*L�@� �g�^ԋ%��9򑪐)���n	4\Um��W��#G��JoW��aH�ԇ��l�o�N��~M?{�$K�Ey�q����'�A�OF�IE�7�'鸲;���N�_�؜W!���F�d�p,��(A˄~�
����2K�H/���bC��/ұ/�9�/�*�`����pOz����bu܊�C�_�I��.��{#?nT��n�4f%�n3�²��B6ٟ���bm���o:�oa��XX�^�t��LO#'�f;������.�W��x���Ȋ���	�� �.U��PL=e�,V+��AC~�h'��h-��L���Y_	V��� �A���.����7��8��P���g���[�HĳNI�M��_�� ����}�S8�o���^&K#>#�	�TԐ��ʮYS�����-7j��ZG�;(M������3+Lv>so�8�
��"Yջ��&��&m��kӖ2�Yr�v@߳圇r 5ց���a����g(ҮD�`V�<`lȲ��|�V�2USP�1�B?#� ���Mc�-�a��][����jpH��0�O��,o��Y����G�	D����K�S)�ͫy".FL�[���\��O�5����?է�Ɂ���5�o�bF�W
K+?f�9% ���C��V8�z��E,��svW!w��O��,��^�~,N�'�pk4y�dJ��K	�t_�]�j-N�m�����kT_�ű����-�C�.K��)��o���CC�͂c�S�zWW�\)�� �Ō����R�W��7��/�uxq���R�����L����f\m_sQu��ȼ:٬w �8i�f���u�b7��D�HDҁ�Y��~�a@ R�6��H����4֣��S�	�8=���#}s�W�}���٪l��h��	?����t�ڈ�GK����v���L7����O�͸�?�`��',Q����qRs�eP��LqN�W
�
��*����Ā�\x�P�8*�4��)��P�Hx�yJ+�@]��}�*� ����sc�һ��'���+��Ǟ��!/r��i��)��.�TG���e/U��Ϟ7 z�!�pL<q��]���'���Ir7ٍ" ����部n�a�J�Z���8�y�a��@�k԰��h!���T�bH�Ș��2��/�#�������S\��*�@|��X�xq��,�TN����k,�`�q,�*N��'�{B+o`�ϗö(�5�������aH$�:��'�%� ���ԕYE����1#� ����:�b���p�N��{�,�Q�t=�T���)��kn�kJ�LW����oBV���΅M%�V �'��7o���c��P�:��L�x9}�[˥�[�w< y�mp���ט���XF�N���f�|F���*��N|*��/��W�y�V�f��-��ZJ�!V{f���̦��O��~��[�\g�^���ٮ���N�2��He���UkZ��9d-3��!�^��q��l�n�&�5�	����)����ˬ���b.!�ǝ}ѹ��� �._�o�<�o�*�z��d��C֊��z���$�����
�r�u�+�u{{8�a�M���<��B�~W�8�I22�Yl�=��g�G���V*]�����X�b�8��O�w�x����eB@�Mm2-��訇<Ā��Pb�}+#b$��ԥ.�Y)������b��6���h��c��q�����*���R�7&l������  �c4�ڌU�/lC�ty��P@5k,E]/'�o��X���n�o�U��$ K��p�ܶ��̘W~�$����A��m�@ⶆ5#�}v��M�u�_!I�o��}�\�ջ!�FZ\�۪m1�p�]�)�E+���oQv�צ?��53`W�)�k�j➈P��|(��s;�A]%I��֟iaȪ�f|=��U�"Ɗ�a�E&L͘��z/bt	�5�Oh�]�QJ�aw�	��H���
�Q>z���U�y���T�c�v��ڏ�Ɖz�k���@�����%s��y]D|Gx~���r��9��9�H��q����(3��(#�=�G�r�I�V���n;U��������H�8��e�g����v�A��t .�g��$�����%��W��[��5!��)K�{;Hx���"��1K�ת�(�` �,A�4��@ќ��C�_z�MNI�/L��"ˌ�E%'nq���h[O]�0;�h�����c�Iݐ��E8U[��
��GP����#��}��؉��g�
G��N��4�&6|l�F"U�σ�'�C�����=�u��j	��/��	>*�a�����c+#5�vm�Ҁ2�A��ggh��ιG��C�K��Ee���cu�k[�G��,"�� r<���i���m]���S��b�k]��Xu׸I�����%�yJ����d�5�� ��_�%}��K2/�)	�#�U�1��� c��=�0;��R{.����y�i�иZ��f3������c�B N7�2�A#�[�=��ϴ%�rw���.$��:g<5x��ߥ�?��D�f&J�k�M��R?��ߛ�m�R8�=��[���.��w@m�lT��YVD��R��}�L��l_X�m㹐�R�s��Ӎ����!Ԥ6~5us)\8��Z? ��5���X�����׷D��k9�*G�eψ�H���h1��5���"[Ο�''�m*���e��
�p}���e�4���&l>%���{��u���x�|�{5K�� �R�,O1Y����2)w;�q�^�ΐ0��Pj��rZh��$�Wg��Ku��>^���vo�7(�g�����*^6lr�}`m���2���m�+GƑ�UD�kgUq���M�<�����[���;�V*��\��+C��A�wp0;pt-{Y��r	�h%${,O{�'B�\� U~����Y�5g���FJ��f��$�K�i���)2�N��*��sb_�)Yj�5�W-�	���\��T�k=����`GO#�72��f �3������˓4��b2���+��wz�e��u;�x:�,���T��G��so���z<���Ծ�p�����7���)�9I.}̓�̀�՗7J�4���֙�0���/-`����0G�rG�n�׏��A��@�#Q���5�Z�
y,�Ϡ�
ԛ�L�a�:��F���f�#;cſ��M�>���a�|����9�1��D0�����5Z{ǆ$��8\n��_�J�˦�_dI�mD--`A�����@����qԍ.e���.1IB���������0D�F�U���]��3]¬S��-6�
��m���׏��s��k�bi
�KiK�&�LB���l���12)'R���"���)�:^�d\Q�mF;tU��{�Wo%yr�$�y�5���<Ϫձ{���R���$Ћ�ƞ�#1��w�Z��`�e��mW���T���I��Ʉ�)��*f�+�.�$F1C�T��b���)����>�@�*��&2e��i���I�	�<.�!O-��4��v2��|oX½�I�S�+���?rm��R[r����m` �����N��Re�BQ_Sr�b��a�'#e�m�GJ���<���fS��kT�%;�0=R�ud�T:U��3��aۤ���1S��}j/��Y�U��H�6�gUCMvj�k��|)��Uy�R\.��ٷWX���12/T��u4E��[¹|�ի�/_�=�!���'�<�+�s���`3</���ś-�%s8�X��4�5e�gU�����ʤ�����-	�7\������Iܼ��R�9�_�[��X��v ?Mo���Gt2��5�R�8����V�^c�#U���
Z4VBM�g�E�Gxם@�A"���zG�9n��ʽ��y�Ǌ,����O����XL]�������ܑ�OȒ�B޽�m�����g�}��Y��26�}Czߍs�U�Lj���r/G�u�	Ҁ��������.\�Z���%�1�����*����7���\xX+��T���m��mq8�A7%�zP)�&]�3�{4C��𰼽�F ���,��.~��90��0�BN<�Pi)��Ĩ�Y02u]@x���K ��%��f�ǥ�'�����䝐�a�ߥ�ӮQ�67f�9dǲ��?�b�m��,&hm�'��5����>��ʣ�)5 4yؙ�[ҟi� _�0�;u��:Ww�t�r�V/k6m�y��N��;'c�(6OE�X��0\�g}�=��z �Z��J=©\��
Ξ��R>j�2Q(�c�u0���'ѩ@z�l:U� a����R���:y�dwd����P<Y�%��J+�a���,�#�u�b[��H����	��[�$���k�y4x��EثXE� ��h_�̇M]Q��	�hm���'o*���� �,�_k�=P�'O���u��
�� ^�S����<���%�r�Hei��|	����� 7|�  ��qh�0Z�8c���)���sl��0�r�3j%N����p���I��LE�EȆ4�®_;��Ӫ���}�w.G�Z��\	��ݭ�������~�1U{������ � J
gq�R��ޣu��p�UVO��N��W� 0��vx�zFj���Ԁf�����w�����<�����e������ɽ�qob�x>Z��u�'�ѯja��m�~^�#}b):�����/�U�#'�Q���uF�,*�e�����;ȳ<JA�X��^W&4aeBZ�K�o`P����M"�ӊ��tA�mo`��,�^��v��ɥ�_O�����cc�Mz�pk�T�G�l#�h����h_j�2�=U��¿�����0�����V�/�d�`h���e`'KU:h��o�_���_�D((�ϾAٔ�ġ�Tg���N�!c��vsǮI�N��z�&�
�Y�+���K�E]�ˣ�̣�=ƍ@ÕG���[q�X��V�o<G]�K����M)J�'k� _�R���T���#V��|�st��v�`מa@ H>��wpw��[+n9�;�o��8�{ވ��N��F�F��[ŀ�h��Rޯ��}yV�B��
�����_�O��;N�m�����d |+-k3�"]рո7H��� }���5Ca��p㬽�Y��o��H+� A��TG�e�OR�����^���0Gx� Z)���2Q4�ܝ��ۍ4]��s����S���EB���]���e(��ס�����	���&zg��d.uǅ�U�����
��Ab	%�\��4�%�����q�u�A@�oS�X�0�u��Բ4�����nt[����Zp���(׌dd_b�����GG_��RM�*�����hgD�w��#���<
7��|�pl���H�H��L��T���7�u�b;Dආ`� t&��x�����#�ץN,[�;/a�P��*�%���-����/ڵ�'�*��7�>�i�>�����>�������^D;fZ����]���.�SJ@fq-3!��d�fOM6���5SP�Ea��� ����c��fn͸-cj+��uN�_"Xy+lB��`�w�5�_�]݂�2w�Ix�T�&������w����4�hׅX�Z�==�0�6X�xT+�	z�3ɻ �E=������O���z<�MxߌC�
]|wSGwK=x�{oo�AmS;+���:5��s7ō���z�x�yH�0��܄��q VAH��ǲ�-T���O!;x�6��o�1�(3�zר����J��ļ���rM��;ɛ8�V��
�,nG=$��qRq]4���`���-���S����B��$��<A����v�[�ܵq��Ǟwb�9Wė�'g����,y||Ub�=�ip�NT����%����[$�9�QJ��b��*�s�`dh�@�)�|*ܸ�}/��,F;����#kQ�[���'���?_�� �m��&�Ӑw��(Lpt�F��^NpY7^t�Q���|\��I��agA��JY<m���7E�"�����.r��Uh�V鎣Dӏ���^����������)��t�� S@9qv`;���'A��A��5\��  �r��0Il���0P��g���N� �O���?���s��UK�����lb�ga���F����i�3�kq��?=1�	�������[�'���@�hB3�-mˍ�{���|6�	Y�<���CQw[!~P�s�9p�UO��Z�m�@��f4�s=��>�]��u�
�qC�X�O����1����9Y������=1�۳��ZUU�2:Z��I����Ko_k��'v�`)��Ǔ�=$#�+r�Ѫ�vqw�~��Sē$\����wW#��ٴLj��`s�dS
����83^�'f�>����?�7bj`�S&��b@��2��j�T�4i�|�B� �캫yo
 ؄l��~�mk^u}2�	�8
�������P&�,F�j<���['�=���պȫ@#297�8�7�㿇���y��q����/������l�q3�1^�hz��o��$��4����߯hb�%;���#{��k	4-K%�M���	��N��t�>E�vvph�������}75ة�:Z�L��[,�hi� ����`H����k$[+!�����W/q+0T��FT��S�4��{)�WcD�+��-ٕQ߈yv87�z�p���`���O)�,�U�.M���o �,���������'�ƺ*P�X� �&�����<������)\)���M��̉�wŝ��F��e�uL��?#\��T��SO���l+���S�$�`"�;-����}�+R���
8�(�Ǎ�u7��Vn?rW@�)2+D�#�����4qS2O����s��ݑ���:i����Tģ���76�P�SAB�*��T�Me�8�u�sUT�,������8�l��U��>71�W�-Ս��J_�r6렔FiA���bDDI����D�'=#8�f�H�R�P5�ufU�B��E�8����b�=p�v!��ksq�����^�sc��I�+wO�z`!=��c��1��di+]t4��0v  ��p�H����Xy�4`� / ���+b�]�kb[�s�5 �1��&|�܇f�7��2��x��_�$N�w�}W�yң��;xD�9�HKrz�S	V/Y���U���C�s�4=R�v஡`Ԋȱ`��W�CWqG����eq:���g��5z��:�
ݷpq�6�C�*�f��7X��G�Uլ��=5�G=����i�:li'����*��K�&]֐�4(�<��[��q4�H�yb�&�6z�)"]u���cCD����ٓ��)�f�����±�^�2 �R��TA͞��]�G����,ࣤ�p�la���i�Qѥ��'1��lY��+��2�rz��"48�s�7��A�Z�UBȔ�����W��kO��qezr�BeT�a������'��B,�	�x�Y����i����I���)t��X��Ɠ��XP�*����7��-a$Lg��������c��܍p7���@����Z����iw�5GVh`5@��j6N�u�O�
c�q`P�ݹ�s�Z��1�p��A��]�j����3LH���jY�i�Ҏ V�}bآ�Z�����div�cB�Ƣ��kj0����~��˄w�s����n�����-c����-���
m-�^������N�^
�J]M����ؠ���:a������Z}����d�.a�*��Д�<å�+�u���J��8���5�$g�=hL[P�G3)� ԭW;$.��Z����QC�WT�0�l��x �V���ֶi�&��٘�=�L������Cv*�;àTDR
��@NK�O�0�����ȝL��zS ���7R<oj֮+��0=e2�WOW��t���Ms}1�WXŀ����#�-C&�_�|C*��/�99�kv�dl�/��8�1��=������4�Q�1���h��6k�e7��7��@��&N�k�����Dec��'���H:��n����X�G^ħz�X�r9�oL���sy�mS w��%ϛ`j<��cA��� W��I+2W�*�J��]�[ k�.�F�oИw�K�S���!�;�G��sR745�¡bv��J��E�L��@�B~I��P�T�.t��:G6�o�<j��L��F�9i�F��B�q����/Tb�ߣ��R>�3ݽ8O�����\0�㙅�����_0�2c�*M���c�i���@S�jh��c���Z0Qq��CK`��$����_�/`R''��^��~SCS�F���؊�a`%�^���#��(q%�uq*rd%�k<� c�_W5$��ߩ�,3��qӟ������@��.$�k��nBR �'%�+���o<�|�\ 4�nɱm~PM^�����У[�<LK��B�R�/<�f0�ZF@�ۧ��n�V�q{G�dv[ ���d4�z�x`�������8������;I��u�#>�[�-�+���j9��.��# V/��S�m���� ޾<n��v�*-/&'���=�G����T>��9�����H�ja���3�����E��S��;u���7��ƻ�O�e�Ԇe�׎�*�M���[�bo�@wS�lm���0џ�mk_����+��}��)����4����_��2�[�ϳ�r`���WW��N�����z���JB�����"��ѤWs��� ��
���@�]�Q��#>	{��,�n�Qg��C.BT�<���'���O+�Z��^o���̝��њ�����>�4x��܌��A���e��J�\�����S-"Ǧ��߱�����r���6���3��K@8���l	>�F�/�Z��r��V\�sI�I��-�QJ\�UݶXI�7����A'y�9r�[�ܿ\�3nY�I��0���S3�NvF�)��R���	�ў��f���N#j^���ٯ�a�$�3a��"l|��	�qU�o �/�12�%�銆�A�p5�p�-h��v�M��\/�)���U�~���A�RROw��x�a$�"O8��8o�-{�mn�el� 0t�
JQ7�y�Ru�FGHQlBaÒ5L'���&3y/����i�A�0���ӊ���cq<ZµT� �����7�/'6�9�2��/e_��;k��+�(R�`h�~�ynY߭����Vum���sb�4����MI�|�ӯ�P]�-��
�h��}DW���hDÇ��VN�Xq��<1�R�T`����-�����.������4U�Ņg�f�%���N�r\IF�q�60����ĝ�$�{-��c=�'��'�B�_~v���\1&{�T�I��^@8���mbj�h��0�R�/`�)���ڨ�}�ބ��������ށB� ��)DQɰԈ�߰vx���
N�$���+� (�ֹ���/��~/�m��@x`W[�_��Rr8��*q\���MS���7[dLp��%zU��zy���49{�Dx��K�����|�J�F��g�Ӓ���k&��jD;�uQV�������.G@��:wt�
G�iѼT`�C;�(#0�t_\^�Bsuc����YF1 �"~�m�>��˅�@�^��x� <2�'h���j�dV��O������>v�=zû��ө?x��O��!�]���J]nIG�kMc�Sp,�֫T�]uD��&^n�bR�3���Y{�W̭�}�aR�!k)�<s/x�w��Vu��U@}���"��[�)L���W�]���j��w�F�=	`e�9�����(�m���{^��CgM���!-�t��r�]˩�>xp�n0=��1
U�|6�8by���M{�&�:p+�2s`O�;��}˄�K����������"@U�B�?����Bz0����r6�`���E�As�!��G�����k���f�L�a��z�,
?>�>ݍ��Lr~4Q�.�̣��䯮���^�
'��Ϭ�O�Cr&a�f�_�e�?�] �2.>��\�|˚�B�\�Mʄ�'�p�l���]���1�|:�C2�#�K|jh]*VCG+�J�0d��e��=#_k�=�V��Y/P���t=�+�p���m'z���?Ƙ�|�\�`�Ao9ɵ�-���礚iij7�)~�`3W�:\��� z���%3��n���yF�bmB���iTqir��J��7fa�� ��N��D�$��'�l�/T331z�Ȩ�϶-.����^d�3�{J�Y˖��J����Me$�v����&����#�!���Cy�" �C��� ใW�(Q3;�O87�rl�P�t?����艛��`\T�+���2�Ȭ��
C�fk'��'�Y[�2"�`?���Q:o߬��X�3E!���j"�݇��V� �á0��&d�5m��*H���)�`|�+%q�5I���PǍ�ƒ�,�`�&yzx����^ _f���nG�J*	w��pm�o����,���ÃP҅Oc$���:l��� �T�EB��a��C�a{v�+ŷ��B]��HqR't�>���<�W\�{�!�z����>R)�{�'�Vz���U9��T[�SԆJ{��1� Odh���'�t�{�`�ԃOrn�%ш��4f�)����N.t}Z��N�ٮ/"Qm��A cҋpz_�����m�EaW N/�#o�^xS������,�ZUR��p̙6y�%"�����nGbY���3�hT�Q�P5�0C<��fB=�9w^�j�D���s�H�Tj.�LCu���E�}F�
�!w����K��BҎ3T��q�+Wα�gn��m/<�h�p��5��9�e�h�������zG-�wE"^F=�i�����O��0
xW�?�,��߿Y-]�Tߞ	H`T�ࣁ~�#�)�/)csګ�T����=�n�y�g,�����_�w9K��G�A��"�l\�ɤ��E޳��[hX�3��[�/SNL���y�m���-�Rjw�5�M�!�m�����q��]�T��
�%��C�ƃW�7V��
����?l�i:v���F�� ٞ5bW��ç@/������,�Y���K���b4;d������J��Yl��ڇ��˩a,���H�7UM�q��c1��0Z��x�Yϯ.�W\(mMX�$�?&��f��z�� �B��F�R�&�1��}E�T���DGPq����J��ĨJ���7.������
|� �X{Ձ`�z���tffR��Jܘm�W�(6��� tO�lw�vҰ�6���_HN�!���\9��/%&H�C����;E9��uc ���@�(������,=&_88E  �����ZZ�<l\�{�ϊ,�
G���f����T�/M�1Cb�[��yR��ɍ�ATr�&=�����^~˖$�N����ɶ�(I8�х3w�]���o@�f���NO�V�`��ŖJ\�㞰^�S��J��F'wA�Y���e͐� ��W$|N�*O9�G���D�"�����/��:rY!(�l�G�1��;�	��Ğ
�EQO_�^>*)T��x ��l�����+gd���x٪cu٩�4Q_x�y������\�-�w27��'�����(���u���,�ժ��c���`�E2Bv�>	��oH�oŨ�����=3'��7�cT�0�"��]j�Y�h�xC�ji��g��ۑ��V��D�1��H�{KM���`����+�,���2.A�.�� )��Q����i��q���va�.�����/V��Qvx7{8�D�3:���c����\��f>��ق+6q����A���GO�d�����yھ�b�P��������ĥ�}��
�Rg���#�ے�� �$�{�ҭ�D*�$yt!��[��ƷP����	!(}��̩),�j�ݪx'��+�KN��c�l�W5�8�����
�xfF,6�;����iz�^<Fw#MlWWT��eFe��Sq�P)����$h7i�]���n�i�8*�n�-��41�0"M�����ْ7�;s��ø����k�Xv��wQ�_ ssS7��+�{���r۞1 ��b�ba�2 ��^�p����Mr3�4���'ݼd���>jb.9|������@��Lg^p�|}���G�Y{g,kQV�j����-M���Jz����Q�P#��n���~�p�$� ����� 9ZDq��4���@��"�&DR��=��pĜ~���*͏��Z�g������=�)�qg#���w�u+M�h�2��\#�@���A�mm���-��v�ʂ	��%5/o�R�><�~+��#U,�=W�����dˣհ|����$!ۇT��	�~[<X6�"|Z�|S� ����(W)�͵����jJ�2]p�C��w��ص�N�mD,��RTM叠��|����K5- *����h?u�q�s��R��y��b����!0I.ε��"�ՓqY�#��g�r��E�!��d��/���1�]��_rs�i���	��Ѓ��=�F�,���}��N��� K�v�+f���:@qt�����n���l��B����#�]$85���?��<\״����i�4�sd$_�����ޝ#�RJ���OL<�)!��_�%�zP���P��Ndĭ�K-�^4X�˛�`�Ņ��vl�39���r�G!�D^����1&�u���~���=����z@�t;L�*��	y�oyw�4��:�E�x�,�Ir9v�Q8

�u�������5}L�#+��כ3��b؋�Z�~�B��8!�P1�G��� ����Cn�Mz�z�K���������e��6�H}?�oW8ox��B�In_Јrϓ� ��\��F��&D_�×0O)��;(SƢNi��a���!Yb��+��G��$l=S	h���磢�s9sI����1�`�%$�n+t�� W\xچ�%W%�F�J��p4�����q�n�W�[���:R{���mWk6l��3Ȳ�%��Ϥ���A���Z!z���� ��Z���AP�wCXc�T_=8G�3�	0f����X�+)B�l�i��ܡ�gR�31� *�����vU<�D)H�����W}���b:����U��Q��(�M�=��.��"E�7x���c��xZCv��4(hO����&F� �GHp�����9���QH��	I��,C	���N�~o�ѶO��~N���x*!��,����ب:����j�R�"t�j4�@Fݫ.o��_�|�#�N9kPӕ�(��K�ei�� 6�`x?��Xo�@`15�lк�?�O��Q�*NZT?苍�)����M�Z��B@�%@ �����:LZf�9��l��w�7���a�f4���::]Z�۴Za�=�	�Gc����)����h-Vǰ���_�A��'��bu��+޻݉n�A�Il4�q|G��
R\_%T�0���q0��ﴈ<���@���{ ��M��L�F�z�YJnB %�P�!�KL#��1ٜ������Y��r��Ǧ���z���]�5Al:-���36b��r�eafG#�g��)�XX���C9v;(�,ê��$��?�p�A�>p�� t4�Ϥ�q��4�B���O9�)�4�e������aE,�Ҧ��9���fA��h�Hq�l~�����ŪpIRWZ+���_�7�����D�Є�^��>����Y_f\�ΡT�o!��
��C�\�� ��[ �ʆLv{{��3ه����'[�˔P�eF���e�|!(�\ڮ�lA��-����~Q(̆��=��>U/�(a�N5��L�m�s���m1�Q��Z�<�;|�iWřS�R	�L�MeI��n�+(�(� �m��1�\�N�<f�@��i�Jz�(e%'�@b&uU���/�  ���{ϟ��߲i}���56kj��0q.~��_��X񲌄��+ĥ��;���|����8�R4ܒ����չ��<nP$�2�z���}.�< PN���o�˕��C�q�%_�O�72I�đ韮d�R�񍿨}���4E4��^���疃YK��/Vg"%)<�h���T��7��=!��u}j�.O�a�v�}�K-�e����O1�����_IE�O�!>øڃb.�]7�v08���X�q�k��4E�$1���h �jU��8:��\�N�,�'E*p��-��M}킼��L�ÁW�c/��%��p�0��������������v�آi?+�`�ܧ_	k�	a��c'�l�"�������н#�o20q��zu9E"+���`�}��W,��]���~DN?���kJ2ϴ���G����_b�R�C��[�[`b�0q��襃�Cb\\���V�h�_��1<�r���S�V��U���}[3�M����`��,��"�[�߿�� �V`v?0����JQCy )��T�w@R�������Rm_Y%V<����:��l��sl���EJ	��8��2��lp�WI]D��ľՉsD���>B�Wl+7>��!QqHH_}CYC�k��f:L�x��4�o+o��Gp����c��uA�#"��\��d��fs��[�_�И���|$�x�����&�E�"���4���{τp��I<NX�A���&�:�A��-fg�&:��$�ȶ���2*�s5MW5����>�?/ɨ��g}�� ��PIĜ�Y{��WW1ф����S!���6+��`я��hL��^=�����}�%���Ǒ���ۘ�XX)��f,�]F*�t�GC=]
�s>�a�T����ݹ�����^�eN�O���M[��
�s�&�yr�Upɳ�O�̖�_fvX�8�~���)�
���^kj�}hŃ�x��E�����]�~�'�dԺ�r��'gP���.@��^j���j`PQ��gJ�8Ky\Q\P��S��r��)i�	t\��ɑO�����S������U�Du���4��e�L�T�\L�ڠ���D����ּ��;��k{��|��-����eҥEH��α� �H��ҕr����	8�c�O���Z4VWy
��9���`���	�L�a�+j[&����O���|C��nI�TV�Md'����<R���M�|�i�Ԗ�	��ɫn��|Ai�{���U,�ê@�?֩/_�=O�3q��A��Bu"���\
��/�@~��o���:��l|��~��W|��vKB(bϖ�҅�5Uk�W�#L��]�1.��uU:0��A����Зa^#��,�9����sO.JX+Y�y��Rb���/hy&�)W\2<�pk�����hy�`4���L���O�VS��?	x�J���j��)���qpжF�:rX�N:oƆ�˖���t]��b��V�xw�8g��cZ�a�4�pU�&� ��j7|��`�ہ�v�-�l��Ƴ@e[z��>��mv��r�*�QW�$&�F�Ǝآ�`�§��p�~��٢jY!�z}\���fd<�! q'���Y�]k�[e;�*M缜J�i��E�9�Y�Ժ}ʔ�Oh�3^m+�C%I���ziw�M�� �5���t�}$	\}ާ3�X��߄����Ulۨ]����e���K/�P�&��D��y���,&�)�+��9W�-Qi�]QbR&�j�4�p|����+���K ��(r��,�/�v���`2���m�zy��鰃�ر��t��^.~�1�� ���U���S�F�������SVG�Z�ũ���L>��)�3����)U��^��%(.�e�K�Z���Yy����2��� xX�Лd�ۈ�D)s͆xA55m&��4ca��X����R�0� ������?���t�ޜ��!��[�k�B|]����e�W�G�ڌr蕒t����!�Z�/��[�I��$�Q�k޾�R�F#��	������d�~u�y9L�|��(�O���aё{��Mx�R�b����4��#h���� �E5Q��#�����y���*~���r��K"\�sq�ϧ�������\����ޣ��:C'��H�N52v�]Z�j�;[�	����w���A���coa(�0.gx�s�+%| �ʥ1I���^�i����[�ǒ�F�|���E,`c��c�NP��{ܯn-7a�7�p��FM����t�B�B��N�D��2��|�u�����!#���=U"_�2F�X��J1�,>�k�����	����&gC�/�k�;V-ѦܱG�� �p��k��
��M:��Aַ�R�B�3�mE�+p���}�!wȄ�g�fl_�;�r=��2��y�m�՚1ZS�*� ����L|W��u��|6�\�����rR���.Z8*�E/gcfLTj��
�����ӏ�ѳi�C+�v�r)�S4Ȥ~�m���b��6\�l��ݝs�w>��W$�]��o�5��1�*-��gELS����1H��.�e�d�ju�ky�W+ʰ{2��67ұ�-kx��iⱄ��ڞD��*��kɁ�>�%�1Y��կ�}�;?6��^��Ϻ�����h���Ҧ_O��Sp���������6�[{zU��=l��.k�C�%�(v�{t���4�����&O=��4r�)���%�n���`�1�p�Zh�E�߸.���}먳V(Mg��c"�I�MP��Y��H�Y���B�
�c� ����G1H��y�lD{E�;��PHY���c�&E����J�f���W�D� <��S̩��|�q�a!�wS��V�x�ڬ|V�/�J�C�Op^�%��_9VY�-��������𵀵�x�� �jЊ�S ����l�����^n/.	����'��f�jQq�#�3����]J]�G�5AK8�b�_�F�{�4�T�S��� K�hYln��y��l`�L���Ԫ�� O�n��#߈n�TV���
�JTܾ��?��W��,H�Q*��{q37�@@ �a$�"X-�W�s|�E2=V�fK���X㎏�.���L�'�Mҭ�Zw��.g�(���j�W�Kڧ�C4�;4�������2���D�Tˊj2D+��f�F� uq�\$wL������ZP�3\�]���H2� T�=T1�
2��V*qc�JP�ܰ@���b�mj��9�v[�f4[g������t=�w�:�!|��DQ����qsщ�|)�_�`Y�	��n��p:�x U;�~=����34�-���k�� 2���_�6l��Xz"-�o�b��"n�b�dl�p���w�5>!=�p�Yqd%?��Ʃ�����W�����P)����A�zhs^Y�M����)L��y�"*sx�1r�,醲�x���]�R�j�b_��m�j]
غ���V���'��<��E���'�&�|��r�,-#�T���*�.�2'��*���B��>��a|$���������>L����Q���g�����uy�-�	�����pb�b_�S�|���繒r>�1�nP{^k�r�S�!�ē���):�f ������E����%�l�3�DB�e��_������, 
~��	�����i��C�Sw2�5�s�����}�#��T��N�ـO6[��q�+��7�-(��a2������@�u��.%*��:�C�鱳F��j�7Q�u�m,���u�\\E�����b�-�>˨��7���P9[���Ex���wEO�OV�����.X�KYL��`�G�R�bd�I=��%=���"�q�Y�	�^��z�;�]�
LN��vi��L�}���G�����^����*�#��`)�c{�ԁ_�SP���t�kz��v%�T"o :��ՅD2c�x��Xx���i��Y}���
��c������>���'����7㸉&�T�F#<u�>� 3V_���Ƥ`�g�q�@~!�H|�����qԴT�����m�'�����}���uW��N]�R����a��u�t��e��]��H��Ne������#��tD$�A�rK0����ڸ{I��ȥk�N��"Ϩ����c���(�p$uG��~*Z �Mv`��+����H����M�����	�1[P�v�����Z3!��e+��l�`
C�,g��h�;8��M��D�4.�p7d��k�T�i����l��~���2Ml�*~�����eɝ�F
G?�(�`Dm�~^��0���Ό�,��"�
����|�����/����J�WEi-�2���ذ������C�H�_|�����֪K�i( ����� @������G���x=��R�53֛��W�C�׼3KV箙��)� ��� i���F��Lκɰ�W�;jbj_R�Q�V�� �y��/�;�Ċ�����b�rU��^��ʤ�I��*��S�@�.�鋐��t�ZAe�Q"��U�mQۏ��k>,j����R���,�ߗ�vy�6�8�bHpt�D�k�����NKV�4�� y��ܲ����.��"�x?��[g��qGT��k_0VNS��w�4P����l[�W)�B171C���h���"���0�gyǠu� ���N�b�a��+���:�6Mx��J��=����/�֦.��7�}VG���X�D���r7���k=M����y��t�3��˃q��6��>�|���*��x!�q��	�̪���0�'����3�)7�h,g_I�?�kp����G��"Q������l�]Ўq*}ֳ	?��> ǡO�������֢I	�ɂA�+�/[!�؍��1�[�h$(�GP��R�4��6�%D:�=�6��sZ��5�:���7Jԛ�<��{#BC���"d_�pr��'\�J)4ę��A�6޼��ΎH	�*m�J���P�h��
��'��TVy%�۷��_�)��HC4���ɺ43�V	;u��Y2t�l�� V�r�����WI�n=� ���Gx�NIfEK:I�%��G�:}zn%��B�/�������-�>t�/29�7F�鞿L��OjLuw
䔋�ҢDXW��;���G���p�:�nE�3�Ն����/�n��}���kD�,:Uڰ:v����0�b�����K8��_����Ĉ%�A�����j�M�������w
{�]�61�b�#Z+���+��0�����@'咓8j�$��%.��Pz�!���h���R{��yT)���N���l_8�����>�m"[��V� ]�ƭFҍ*�>2����t���@�o(R;��׹�O���8�\]͊(��q�
���T5���,]����_nY�u}rH��u=ʰ%�n�V��Ծ���ׁ�{�s<n.�%���s��=ǋ�+��H3>J��v�����k��B����,��K��E�q���v�w���w���M$d�����6n2aD��*Ԋ5J?��:k�m!��ִa첋�c�e��eb�M�pi4q(�zA����N���l~�Xo�q�]�;#�}c$Ŕ*,�d���jP�fM@����/�q��B��;�R��S�E�tzf0^�p3�e��WU4�	L�Ss4��J���)S̎<
����ǀ�+�����{��|^�p���}޾�N�����"K�������<U���-����ZW��Y�� �P*�M%m���#9/��$9�3�E6!b�Pb�������Hi��!V�Y����V����L�]fB�p7�&�1R�&cSed����*}�] 0ߺ:��dӺ���f]�.�rƬ;F����_��!!l� S�2]���F= R�WR��3�saf�W�SyB?h���h���p�T�Ϋ���m�6~p��� Op�ʗ(����_S��~*
k1ʃ�������mi��v�XY���h�$����H`v�B	�����E�w��i`��T%g���$Dv`o&:�y��U*?Օ�h}���r���WNv���lAx��E���bxh�%����4�C}OZۿ4��B�qȰ �ǿX�ii�g��f����t�I��G��h
El���qC��~�K���(�z�*��PJ�L��������I}�*�@�*�����
߶oP� �:�r�[p�~)�DH�/x'Y`#3O�492
��cn��oT��	m����g=�{�>�s��./�9�t�܄��{���;�G�/�4�|'<|�������^7�	P�=�f�D�m2NG�^�`
�Mu��6^I.��V�ƿL����@.��L?���D�il�&��'~��nR ���h9�x��l�(E����0<s��b_��.K GI�l�L2u/�&�j�qx2`����e��O\��8���b
,B?{=G]��|�1���)O��.V���c��2%�
���S�w�&���QZ���A�@�hV(��>�G��w�����zf~�����<x�m�����5_���6JQ��=�(����c�h����\�B�g.���	�9��a���A>4�5��v�6�R�2�P�*OO�qϵ�ͻW0c��[,�I�濾52�q����k�N�	iv�ȭ�I�ܓ�jf���S�GN�vNT���擬�N&�MږC���1�.��-�ޝ��YxM&�v�#y���ʵ6� ����BV�l�4�@���Ū���S�S�j�7��,)V�{��ғ ����׀��	�25:g�c_����?e��?X���Ogt]�O�s�Q�I��G�qz�WF@���\
�xB��-���i�.�߾���Q�� /3�t��,Cq��Z�qؔ ��8φ�)	�c���^R6|0m�"~Mc2;��G�@H�}^�+�x��ʷ�zi�
V�h�!MjT4�����Na39-6g�y9~Z~��$ls��m����d4�9z�h:�: ��Jt�z��&�NRo��|��1+��K���>�PXQܷ����N[��j������Y����ܺ���U�i���(̈́Võ�Pv$���P�tS����.s��'(�~q��"�����sK��K`moC�X��8��+�0��?��<�S���f�@�lD�T�U3#��!����K�E��B
hk����M7^�ϗC]Y�]V�=1~l�\�c�������E�6�8kH?�J�C��WT���U�)��)�ޯ�y�N�c�bY��[�qd ����ȓ������Uu�Qf����c@9]?q#�ܻ$�����k�����^�ƂCP�RШeC ��E���:���F�*ImM��\��_V��:�D#uRH��$�Ȱ?��-iGC�>�]E�q4Nm\ш+�C��79���ޗ�5���q#���֑��_��{�ɼ	�3\T0`�p���^�ه9�~�'�U�}�u��ƀsPjA�p��SdR X��ÐKۚ�R�+8��	f������"v��#! ��pM���%��u����y��i3�\�|��z�+(L�
ȹ��ܺd�P C~V%i���+
 ��5���Cw5��i�v�mGfg|����9A��1
0�S�h7I�����c����6���8&��c��V�b�~ں��R�70Q��ݸ&�7��R�Ǘؕ2Qnm��RWc�'Κ`�1����	%��~\W*1������� U�Mؑ����il�Gt���ӤY�	�oCU��OdA/i-����<�i�j����9W�u����j����Ě�}.�,a�{�}�$gANok�(s�%�vY�#I�@�w[E�eT�l�w�L"�69�v�Y�ssE�=�UfW����@1mw|[t��.��?�3�I���MZ0��n}{"6J���tc1�ۆ⮚尗*".��[��u�I����{����U:�ݎVeka���j�d�eüx�vD �|�=l�"7��`�8���㱱f�{	�f�hy9.�2�:��+��a���%��H8j4��ԅ�b��URr��;����}w�P߇�t��mC_:]7��q0ċכ;��bA�5��ua��M�[��˦��P×Z�8Z@�W
bք�6���z����_akiz-'�����O �K��*��+E�/ �a�T��������Ett�y)'��+�����ȣ�ޭ��gI� ��h)Il�{��+b���Y��^�;�`��p/ec�+#k~e�/�
���P��A*p��$��űevT��Xz��U9[��2Ø��<?���Xw��gQ���B�[eR��c/Ml����K��AYA�qf��H���U vJ+,q��np���sDoT*3A9(��ٱ'�W����u^W�yŉ��jо��C~9T ���&6�'�y����D���w~�WR9ǃ�Wd�޹R����\���r�������s#�I�eX��;$��'��U�g�
��{	��%����-�oR��-�=�2+����6Ŕ0�f���5�&���o�N�&=$��kj��K��qHMjԈ����v*��E��� ���B��J���8�4>н�X�r�4��1�t�xi"�[����'���H�Zꔯ�62��}�B�[��c�K�(�^89`�6 �Z��g��L衢�ê���?%UIZ�BZH�A?���)ҏt��a�sۆ0��g:1YV���<0�R��x�xGp����f*�;�":��9 �T�Z�nc^¦���q	���AS?^ڑޥL�0r+����4"=����+WX�Sn�ٴ��t�qv���6��G�A�Ҟ7Pe�6��ņ-.=g�Th�۾��S�QIm���C8�?�𪲳��|��YU�2���ڃ���+g�%��;R�tr ,/G�(MB���>ݟ�_��\uM(�n
�G
�0y������O ��k���¶�X�s��Ǧ���n�`��z�E@�EZ7�R�SJ��tL�x�u��ߓ�X�u&�0Г�},D38Q��H[�^��$�p������<r�?fέw�[�l�5?���6������AA.���W�����yK�|�_3�DTs�X,�6�ķ%�&^�:LB�Vc�1����"�n�@��6h�Z���pfU�v�>G���\y6�e����������k��0����|��ô�t(\��WYQ���\���!���L俆F�r�j|^�S�ZO��$��v�i}	H�>�t\�uqy!BD��&�:��X�A�4�qf�4
�-�Yx�r�nA%!���k��C�6J�v�?�u5�"<rD��v_}sW�Fk�f}�U�����u0p?U�:ـ��-*{+7\��;�OHWр�dRym4��2>ă��G���6���v;�[� �>>�����qOz���mD�Y�/��Lvҥ�y�1@�?b�;['����^�ǿ5���k�eۅ@�9��Tr��1��%#�l�O���Q�w���Où�[����M���ſ�}H����������0�I�'<��u�D�ɋ����͉'���1DE�`��^,���%�L�J~R�v��S���q�g�X�����<�u��eH�H��_N�wI&>�iܷF���]��̓��Gd'�b~.��5�&Ǩk����NC��"�M���)+E�iĘ�QA��t"���j8����ҩ��r:K ��3�K��������b�̧�Г�&��]�|���Q��$��\�F����Ȭ����:}y��¢�>l}� $��d)�����iz�)��U<]q��\�kb3Ǵ����f9.�m��oH��x)tݛ��z<x�����H,rS��y����:�0y3�ǝg�31�e���Go|8�ʝ�>H�v���@7��p�ؕ�E�Gv�AѦ��p�O*<RDW%pB���!g?,��3����辎0^oT��ũV���k�ҫ[��^"�^�ZVX�r���
/����K#��O˭�݆eBU׶�7ؕ�p	X�z�u��>������T6=�^2�O��{v����8�F��@�S��-:���r��V ��~�K�����>��F��E�O�GOt�\��;Tj���T��k=�'[�s�g�W�$�AR��Ą��G�΄W�Z�����=����#�e��&��!|����KM�pN���<��9L[u��?��E���̖�S�e��u�j�þgQ(L/�r��U�d�}�9�1oW�5�~'�b�n��tu�-�!��OW��ȼ��n�H��0n�ݟ�8L?�1U����C14t����@�Qd)��B7-���g'AR�_n���W<J�C-�9��H���v�V�ݴY�/U�^2�X�rD	������c�nM�{+�(� ��=��£��5}*}FyK��O���`I㺓�<L;h�u����nh����Өb��88M:z�L�آF��tʏ�a���n�R�8c�y�ߒ�6b�DcJvlh@X�k� ��;�a@#�h����(����Uq�0�)8��J�|��9}���d�������F.Pl<_���Q��(�ߦpE*i>���[�e��y5��H3c��^�봒�e�<Po�+w�3�O��<�C�AP�j�Drt>_^���ȕP���UBĕ�\Z��7#��D�d��B{԰���Y6��|E`������\���=y�kޜ�4���%����R����ʚ���Z���"g<[ aF�%a�V-p��v�O|Ƙ/!�~IY,��|h�ƒFy�£Ϳ�HQ��b������5��ج�fxLճ�{y��*(��&���, i����h6\l������N����Zb!Ώ� �/�*|���l�5�o"��?I>�}�h �����[��9���W�ĕ~�,f�=��+���{��^c8��X?���aTP�t�5������?8�w�O����be��~a�z$?7�A5��m;u&8N������F� q��8�I_$�+p�������'�欑J��
�4�\ۂ��kM����P����Pݩ�+���F3�a1;5����즜L��<ٛ�b�߀3�e$q��e��A����%A5�Zy���GR$Vu�1@$ �����z��$	o��`�g�����=������m����y�6�-��R�zO��g�	�	R��D����'�3�b�~�
�aWt�!>4�f��q��[
��!u^@y�\hc�}M�����U������˫#Y�K��}8��a������^�x�o�.��K�ڴ+��M�'�Vi��Ypn���X�s�*�&�=Ĕ���~>rl���u(	���Ƙ�i�#��7��@��x��G����а5��QZ_%ɑ����?et"��t����[�W�!Z﨑�|'aR�6'��OD�F�S�� 5z�S����	�N��닯�ᑮ���mG3��	�M��e��{h,��32z�	QAv��g���_�
l#����e'(��X�#d�g�R�$�I��z�o8L)\����Q<?�6�P5�*�]c����.��:����U^%浮g?{Dɢ��2L+]�h��	P�ăi��pɓ�2����d	�� ����*��?��f�C��L��κ=@�%y!oG�A}d�2d+����e� ���J�dŴ'����cH
�_�i�~p�-���T�|l>{-�I��7�{h��*������g}��-JA��M�3)���3���x�@↟��b뗣C�@�B�����#	g� S��3��Z�	O���6r�eï�s��2�o�]ܣWB�� V����<������b�12�b����`��7eM�_|ys3�b���w\{�ww��OG�F�H��F%3v��d�A��hQ��h$Zkw�W���z��Tw6G����a�Bսisҍ�8Y؏� ^�-��e����<��m{#�@(���刻nNDqS�D���u3W����3>��^ކ�ɏ8=H<�����մ���s#j]Gb~����X}/��|�$I'�j��0�oj풠 &3O#r��OUgf�,�a<r�R��$�	���ʞ�1�5�X��oA �%���M��ܙFO*[��u��҆/�Tv)���x&;�$����{�.�)qY��4Y2("��!d����f9&�͑��}�9�)Ϯʢ��_��5�4��e���i {��`$�
�-�1j
wn�]�O�0p��j��@�/�*���A�� ��J59!�q
�%?��jzc��9���_�(�e~�75j���+c{d�Vl���L�;*�*�@$	�-m�ժT��=��˲zE
�\o&�6���Y�X:\A��G�Y(-zj}l�$��UHz[Y�yp~zwM�j-+ˬ? �
��8���.l�_q)Lk��n�]�7I�Cp�S-�����Z����#]�#S�u�1%�f���Ⱦ#�E��m0��s6*
�F�k�)sFļ�S"2�664v�ՙ�yѠf=�d�A��#7�Ҋd�[���"�-]P���f�>�t�n�	/��jG����tYvf8��6qX�8pMg�*+I��w}��#��Y�L�`�N��qʷ�t���u=�Vܨ��g�;������,,�U��)-M�3d�%���0�a'�Q�A�Q%h����Yd.8A����;L��du���v��S4n���ӝ�)i�۴2�F�?a)���aD�W��}j)�$�-�s/JI���͎�;��7��k������b�fo��K@P�w�������LZ�z��;�`:�L�{|8��-���P���SM}�:��a*b���i�>E �'bos��y�2�]� 0�Q�ӥLD�j`�b۠�b�8M5U,�t?tV���Y��C_�[����!+��J&)Oͦ��~x�~�������� L�J^��=��M�廊��i����N��^`��V-Pʧ�g�>d�H)���o�^�i5�ptC���lib���[_�$a
�}F�ڀ�^b.����-��õ����!�oJy<�m�� �e8gP�6��yrH1���!�|�Eм���AR-���@�[�5��|���Ҟ]ә�V8ExhRk�y7���ui�'�� �-�	]���q��@}���I���\z�Nf8�<��$B�k����	K��&��63.����?��8��\�*\��Z51>��$�t���%�k������I�x�w���G�0D�M(�T�p��W&�����&u�C���=��/E�V]��u�R�rA� �ߜ��
���G�l���d��W�k�r%��1�îZ���H����x�N�u
��Z���lB�OƬ�
���j�W��#L�W����E�uS��&�ee�](j��y({�(i~@$�)��^���u�DQ����9:|2,{v����lq�6孂i�L}��vb{��C����u��|jI�����&H��\e�\�h&j�JjB���#�.ԺHWщ�D�*58�roG����{@���3GOA���z�*��F#��Ex��9��YF���3`÷7�綏G���EI'k9��W��M�z��Z�o�v`:0I$���t��2V�t	� ��eՒj�Q��W:�V_*�y�������X��Oը�|����2o�&�,x��p$+�y?Ò��W�vR�M�$����Ӳ|���۵��
�D�j���nŽ_w.Z�9��㎎�eKB�$ә�y�x����3Shؼ��_�LX8���;˦`@��ZK�$Of>�j��l#�����X+���:�V��]�m�n��/N��ن���C��՝�m�iK>��>i8�~&I�8���
��(ezBv�6TE�F��al&3$��_�"u�/�=H���@�v����o��}�h�ۈ���ZcE��jջ)@��=p��FC
�X-�!B�Z,+�ˬE�G��k	��kJ+m�����u&@�M�:&�@4�RUwu�Ho=�0X�N	��������=K��M�����/c�C�g�j��8�.�ۏn�0�j+���3��(B�$��^�(�����_��K�q>D����h� 2���1���_�3�>��F�4|��f:��� O2@��Cf;�|7J���	�k����W�\�"2}m<����3t�z�%��9��m�Ti� U6e�32�!���g�נ[t �r�-Ȓ�϶��g���\��$u�-�Bm���� ����~�h-鳵M���2PI�E�df�����.�i�@fV_����]���\:�n�{��G�oz��0�⯏���P�(i ���϶�9F:�FԾYҮ��w_��S� �R�� js�c��j���ļ�f���_(/(�63j� FJ�cۧd���b21D�YClr�f���}� .,5n��v;�V�ms'��X���<�*eu'H�̬e�K�lK8*)~kw#ֆS���G�
/f���˸�,ꉙFlCpܶj�1�)VSf7���e�t-�3�.GZf��>/�c��u�8�Y1�r	wGZ�\e�e_��J;�g�tTA�_��z�P`r��5t�
�e&�|��vJ��ܲ�$�o(ڮF� �5��]�E+���/	�U����N���i5!?�m=��9�M��9'e��Y@���7u�ྭ��ɛe�G��i���5D�	�%�}���]`\q�CX�o��� ��*����ӓ�?eb6t�hÚ��v�8QV^X�2�$����q�_������wM Œ^�Q�<>rg��!�S7M��.|��)�=D�i�CP(t�?��Ь��ʖ����VM���S��qɅ���u��QUJ���V��۰����ܿ����>�Z׿t���\���q�z���ѫc�ٰmņ0hhn���Ѻ�~o�76�^.K�">��d�FʾGhS�w�;�(ZfV���̬P�Pz���뻜��]��˥7�}�qq����:9<�צY��Y�|b��@���u�$���UJ>I&YSFJP���m
Zk8��g�P=R�&�+��p�Z$�KO݊t����lŀG�hgY��V|��f�Kr����Ud��?����շL� �A�1�+H�S,�*����TWƈA��<���Vn�Y#��L`����&�)=jN|3�H�G`�4�b%�ϩ�9���7�ij����8ʸ����ʰ�I:>\���l/Qox��`���З�Iq�`*�����m�}�^掰f�]P���׺$�{A͇�$��j9o,�����҂��D��n�PnjF\W-�Y񫪷�nX�g�ld�����SӐa?�l�ׂc'����F��<tH����[�Z��h�?�8r�]���t�ۮ��g��)��QH�_�g�ĿuH��7B%������Y�J�D����N��ɠ�Q>�T�4������#�"D�u&��_׉�So�g+�R�x��ڹ���������UH�@IB�#�0]-dO2�~�K�|� �Jd$�Z)^�2�XԐ�;��b���o�(��S�ZT���,�C�a�=�-$�����=� �Sxy�;8�:��,^��oZ$P�>�=���j<�Q�6f$[@k���K v�����NS׼%'�SZbg���qֲ|���U�\T\I:�vR�9�%��W@��W��v<ݽ%<�6�&��M*��}�V�=z��o�"P��
�:W"3��c~�z�ϥ��q��ogQʣ���xTDW��V����+���(�
�Br��`=!�����GA:�QF�'�l�=l+cJ�sqI� {��2�(%L<ͩ(���>�b�g��#�V��h�3m���-+�A�GJ�I�L��c�<�~Kʭ�=a�(z��e%j��F)/b4p<;��:��to(9Z(�	ևZ+�6��+���+L)\��Z\����	>��# �*{�,}N@�?���G�Ė����JOʒ�X1z�I5�����W(����-�k�W��}�m�dz"U~�3ǸIY�F�x��d0��0)!�l�g�����(�|f}�<�,O�ѳ�kv��<N�����#^�2�;-��-U0&q��m{'�:����1�4v�ߠ� Ȃ8����*� ����k����	w('�]A�[e��t\�ш9$����ʬ!_����7��&~��U�nYG�L�j���5�t�t}t�e\���F��,��"w�b4SJ"o�44j��������#�+Q�C �9�d< ���첿i�Ҟ�6Z9YN-HԦ�<�o�R��q�o��10��	���ӠG�8�I,K�`=�#`�ķ;�؂ӎ��n���NM�Tڠ��g��G�i�Lx�c�4U���^f!:��8=��?J~`+�!�,��c��.B�+��d� ��f�̦�KBZ 6U��5qJ�:�uaa�Nak<�����Y;4 �H焸�ϊ�*�#���iǧ8񌀮��I)��Ϫ���!;�mr�Km�T�8����<��w�L�
���.�k��d9�4���}�E��߸�u�zL28T�5Rz�R�`�o
�!F뿟9��&j�x
U����yZ�+���x��`��"��f��@�8�i7��UxTq(',V���H/���H��=�u�nN��`gS_�>�ؿB{+�|�=���]������U�~*����
fT�Ci��h��(U!���<�w2�"��Y����Rs�z��j���P�RP�;�Ri�iCr�ÎI0n���۴�I"ꄉtC��E��؊r�.�<NW�εF��V��d7�x���K�a�V�Γ>����ة�Yx�z^UħP}U���M� 1JNX���I�#����w�	r�!���V�ib�؊�	��c�S)�)����jS�4�K���׋d[G��<ӯ�\�+��=q���0^,
؛���"�i� �s�R�f:��`Q�̒d�%���\ 3��V����Ccd���2�eڂ���y;��q֌
�	Rޖ�hx���O�nB�Iz*E�!~^��tj0Hl�Ro�S|Q<+-(	���0U�VU�����@����>zd��0���4sp*̬�����Z�E1eX��フY|���������1�����ɪ��J�ڨ����������ʷ*7���p��t��b�,I�V�,i���X2 �G��c�J�-x+�=N�.!T�WC�*[�����c����<�>��@��(�_ԣ���8HRSɱP��=���@�<��߆iR���������烍lF��fs�j� q����e���fy�����	q�5?=�7Sh�B#�4�1�����E�G��
e��YpW���A��;�����3	Q<���S��,g��G�'syAgc���Yd�%�ѕ�ڻP�~�X/���)� ����Ͳ��d77�4���a�zW9ȿ���4�r� �ėRC�,*���ŀUw���B���)n�j]�kJ�����F�m˕���;P[��5)�� �g���{D
0�~��7����%p�j���iθ����֜[m"A8�0��R��n�Y��(k1����Zr�ft��g�|�iV�����ڭx�����:��m���+͎��z>3.�C��R��|�9c:�A�A*7�uF~?���r�Q�E��p���+�z e��#��6PW�%<ځR<�#�ќw���{S���{��r�����[%>(~��x�Z�/��="��|$�B'ec��4���N�ӣv`-��#���->�=މ�Z=C"I�Ӌ��!s�.`�3�[`54�1�a�(*�(߹�2�[� *Ig�v*�R�?b)�Dd��I���/T�9��10�D`d�G���w5�4��$՝۴P$�}���*�\�b�U�[�Tt���x����?���x������Wd"����q��2HܷI.f�5Y�Вd(/��z��9��
<��'n1GMH���8sH`=���mdaZ��S�)O��e;�����dt��IY4��T�A�x��/�>S�;y�#TG�4ρڈ[;/�6F������fT%@\��N�ew�� `�0gD�x�.�2Y,����S#�5�5mk�`�[��Y�)v�$_?݅�c���%�iZx\��n����{�SG��xR�նL=�Z��Ic�c���sz�8��c`�%��4]���o2ra;�LfAg���y�L"���O0�w�=��|?`�ޱ��c�׃����Ļ�a^��&��Y1j�p��u�'l��gq� �Rp�?�|�[͸m
7b�'����O:BN�ԇBe���_ɸ��=��ti�ԏ�(��~~_���v�vh��Ni��r�˵Msc���>�Ϫm��#��"G�%���%M9 n����fy��?Ѽz�	 ����	�c����!,i�|�R�}j!�3X|8^ۄ��.?L�Z�y�;<K�l� ���f�*��0�U�(���_�\�Q�u6ʂxk�Q�SC��gC�T�|`Rٖ�"�1��Fӫ����My��S4̖�E4E� �v�<rA-��0g�JB��n��;j8M��z�',_�xbM�./O���	ޡ+,6����R����j��������k�C"q����f�U���P1�{r/bi��c�_\x�=O_�����-��F,��.�w����F9��R�!c�Fl�󹬶y����	]Ul]�g�;S�;D?P�O�����26d��FT�.�r ϡ�6�F����|:7�z	��7��g��;eq�⒒�r6�OENHm�^�w�Ȣ��L�d�������F�뿀��;������$h3������%�Ę���h[�����j [wn�e���]F'.T{���_$1,��y �5�@~򍬍�ˌ_�?C�G^����)�ۅR�����"�K�p������[ԉW�o�Ķ�ߟ+^�yc���S.0*��|�Չ�9 f���SWK�g0����!O!�%�s-�M�h�&d��������̠i=f]U�u�͖E�B��J��U�\������ϓ3��OE����Bbc��8�6� ��cyU}h5L��{�9,�ܦ����X��21�/�H$=0f�T��^~i��<
'�
q�\,��HNy��q+���qw�:����%�2��Q�m�O�����(�Ϣ�4��c ��=(�a�ȳ�tN/f�ٳ������H�gݎ�F��l��~�����6�Lo�L�@���Õ&����;����3h@��]�Q�.R�?
9�Z'�8z.V UlK�DƹO�R���3��!�}��Dj����	9*l�y"M�u9v��oo�THie8	��\�us��	�Л:"1q�n�� )m��E�l7W�Xz0�0���[{1Z%lԫ�]աѴ����8��T��I>P����^�Q"�_���!RΤ��ݯ��_�:�bѷD�5L���2ڞ�'�_��CB��+�6w+X3�-.�!�ݓ�/�(m;����܆��ޟ�!l5�l����ݬ�S��8���L�f2?Tw��HAc������+�
�ڼ�Dy��q��.�Qq��C�e~��C��S��L�yU~���B�R��6����#%�m,</7U��9�a���h�$[���w�
b�.�N�]����@$��$���WiR���@_
�X?��}5�^����%��QH�D��疭뎩nR����V~|6P��t&��w��~����a����tg|N.��R����جaViMx�611��rF�4�)���os�XB���L��JC������(l%ߧ7VV�\	G��o���~�G����������HE����ƚ&�	y�Q�j��A]q���Ѭ����T\��j8�������'{;?��:��8#��tEf�j�E���+$"��580����g��*\�d�V&��'�w�dtZ�����ɭJ#�w/���Vj����a\t p�����M�H� ���Hx���
��rEA${��kV2�$�٫�S��+J�[�s==(O?xUu����/ab��K�/m��pب�J���O���;��ӊgk�x_\Ϭ]�:��! Ȁ�$��r�y����R̜�1h��>DY��tI�E ����z]A��Tɻy���Ma��/��*�U�˴�ԛ0F�$#2N�(�ؠ��Ѹ�>
B�Y�+�%D��zT��42��m�ڮ�� �&-Y�J%jYhZ�Q��W*�
��xQ�z���4���8�}��!b���E2ޫ�ԉ3���Z�R��[x�y`iY�OGrd7������u·�~s:�Ճ�Q4~��LD�g��F8�zQ(Fb-y�������v�����$gި�k�����X�a�vJ����Zi�k_�u��r�F2a�y�#ȼ��#׵Th��C^t9��#d.��]�.�Z M�"�Z����d뚋�o�|�ETR�yk�u������2����6X�7k�!���u��Q䜄��p�o�}��Q6��aq9��<��~�7�ɛ"����:���Ԩ������,�,�x9��t>���C��B	���;�i�/�8�V�n�{4��
�%�.	j�E��ٞ�O!'֮K<V��Ϥ}�\�U�3"��
a��f�8�bH��f��S�-�{��ʷ|��Y��Q�&��h�T�eX��0���7}^�^��\�:�|���� �� Q�k��N
�_t����cMl� �zָ�!�okXi�BT6|�NVw�@@5��za�{�@�;�i<E޲_ւW-HCA)Ĵ��<�����yMp���Hb;��˽9Dr��>�:2�M�DPh;8��}�S��7 p�8�3X�?��� ��1�������!~d�����PZ���-�'���p:��Քu����v"��nV��@�4l%��Β�N�硪ޞ%N��E����\c���i�*(�,�q���j�T;��!�6��!�t,��{�ŗj���}R�J�I�IM�3�b�:��x�������.���K�*����^c  �6rj#�8�Y�	R5qW�����(0/����GDq���_�lVF'
�nk�!��
&Y�@�j?�`�{��7jҲzӲ\z���`�����_hnW�b�%5\3�9�l�k���ݢ`gΙ�0E�>g����~���ب���^8�/�K���j5YȬ ډ��z����U+�I'U��u���@Vq7�~:�~]L����Ə���KYU@W��*.��5l@��I�r��2j�{{������B��/Z�KH�����-J�Q�/'�����X���^�bp<��W��Y��_B�w�<�U�>��M��r�}�f|����}�a����9D�SzG�iK��0�o�Ɯ#�!훵`m�І�5���O*�����O��C�ϊ���b�#w`>/�;��_ {u����u����.Tr����Ûw�rm�X��h�djY5��!{x�`�rk���d�
�����V|\Vމ7j�҄�Q��oֻ�B�����d,��X�9D?)#̍�`oP<.��M7�Ԇ(���d%M�.��a�͐Uŝ�L:u��|w��zi�ۆD�ض�5���k��ӳ�&.�f7����V���z�5�XU+�|عJ�7��g)/j(�@Ľ��?
����ʆ"K9��� �����U�y�	3yL5�1�[?��u`f�H/����`�}Vf��%+���N��DVe_A�a�uuB���	md�?�u��Z�6S?߱�Y}�Dr�ѡ�>���o�#���c���v	7w��si-E�87%�w%t弽�|��<�F��/���R��auk�� �Si׉����杀eHX.����np)�b�x�5;�W�)p5�\�XG�h�@І��j<ҍ�x�>�Chx�,�:�og/ܨ/'�Ǖ6/�M�_���Ԃ�uW��]B�o\"&�͓r^{������[�&���W���<���q���� �y�.�b.T�3�D T~�9X��y�T����%�M����3�\M���E�#
�<��Lbv+^��Wϼ�[e�������_�X�d3�I��8�g����9j�M�"W�O��駓{ׄ%+T&�^P@���L�7�ՊЋA�\�|0S���@�(�gN-���M�<��8����j8,{��U���z���z�n`Hn;�-?σ�쐈����^a�Q f'p���:T�d��p��k؎6��]���:�Z�G�3BȑeDeϽt�s	(��פ��9I���������>�+Ąw}�uu������9�O�ƶ�"Sk۾���cz����(ަ�ՠ��n~��S��������l�c>���E����y�a���$ C��A�$��x�'F'㹇}9�Q�A �H�k֣����S������2�/9�����ͅ�w��%��W���Z���^�/M��Y�(�
��?�kI�����@��Òΐ��,(��9"��HΆ�_S��r<hQ{ ���g��a��2+H�9`��@�Qp�m���h2��O�+��I�t�::ޖ3��J%��Y6qY��G��9J��J��WBb��a��
��2ָ1-�����]f�ȖS�V���=!�:���J��`E7>����� Jo�`a���2�6i�q��
Z�������9/��L�]�=BA6cfm�� ~���k������y��E4��}�o�6����FE�$��ʷ��v�Td�kٰ� j�+���
h��BS~���_�旧up�{��{l�l���8Tq�<���5� ��k? y���U��O�rm򓼇@�$��̀)�:���9*e�5Y�u?	9�y��Y:ʫ�I�˻����f�xY.E�.�\(N�[cZ���E��]?�S_��\MB�w�d�-�9���s�Q�>m+�̙�e�^L�덛m���P:��Re�0�<x����v~7��q��W��!BW+k*F�p��Ƶ9�Tel�*�Hx�w��sU���B�m�"�J#�썗y���������{�Y?46��
C�gnO��T�*b�W$�j(PFѵ
��3�P ����9@r0X����Q��w���"$�����{��+C}��a��׻�|�	��4�JF��h+"��f�>�������o��f[9��6���B���ؼt9��N�Ӫ�)� �|go����3�*a���I�i�9����#YI�l
�1���?������&�o�6��	T pڦ%�c(�q��k��<Aз�yK���:t��4�Ȇ��T�cȓ��_2�)e�4�D���3�K.a5t]���l�M=sЈ�l����~&��}�}�-��O�cE\�4c��R���4q�Rގ¦�p?��0����p~�Xf��'�5�R̭����U���8Yk�ʤ�T����~l��4顣~��g���~;�1;�T�^������QO���so&e���Nf(�䘨w��T˽
"�=������͙hq�W��a�_N%���^f�:�~_�\���%J�e�R���\�V�(41n���wI`���݃����2�+�N^V���T�H�E�o���������P�����e?6�����,��Fā�+��H�gQc�2��^:٬����>4C�Od��*<�,�;ߞԬ�rC�~$���|{���3T,̑�r���S��G��Ʃr��纤�=2nn)���%E=P���h�Mʷ���v�[����,�ƫ2�����)hMS�y���|�#	����m���U�?p�er�:;�Q��fֺO�j`3G�"D=oA*f%��*G�?w<�LF��3�Mk��?F�f�|��3$Vz��O�W9���~�p5B����X�8+��տa' A]��q��%B���LU�^ʛ�\�S����l��w
�*���.1k�ϔ��� �R�� 3�P��!���+�s��7�So[�d��ԇ�����;�hK��ة(H��x4H,`��L	� �s�(�<�[�^���_�R*��v��BP
�}cyʗ%S�b���}(��(�c�%���{�$-�m�S]�E:�\:l�][��(�617l���2�xƄ#Q'�gϛ�$�9V���+���>�9{��Z��n٘ƭ�\�s$��ķӑ�g�p�Q����in>�2�S�+��\�9l�\�1k�_.�F�w��䎝���%~J}���������qRN�f���^==,��qv�ٰ�c�I�Y �loW�Zޭ����RI�lq��#�+�ǲ>���4�C#$dT�;�Ӟ�P�eZIeq��[�|_5�������Z�UY��\�e���V�6���~��J\���'�����[��:���˭w�,_�j�`V�W 0��l%�-��ܫ�4�ɫ�d��.�.[��m?w��F"*驥�UZhĬt�/ A�f�V)�5�I�GF�3�^C1!r�S��F�P�]V��#��u�ǈ���C'LJŭ�Đ�-'�J[��(5�����}���	VDt�5ױ����[��1�|Z!(TV��4�ん���k����#&
q�휋��sIeg�iV��8`	r�6��i���{�&���<�����.o����5~dKN
	kj]si�M*A�ʓ�:�����Q�3���Z	b�Y��k�9Y���
`Q6���"p\a$g(;�Zq1[����RHx���4�n܊YJ#��R��u���k���Ce�Е����NP���or��R�z�JI��W��ה��������I��e&i��HNQ�jnssk����Q'!���hjq��?Vr����	��O�%��|E��#?ڍ���9Ī�a��M�b:Rt�Mm��A��u�G�5�7՟�'� �ߛ*R�����.�> ���V����C��m=*J,�ִ����ЈA�9����V�"��ӂ���O��}
YH�)�P^o66��]�Nm���2w�@�(%tID*J*� ���5!~?l��Agf���Awp�e���x'��F]�U�Q3�k������X��M�:%�|�(�>��Ղ���㎎���3��!I��`8W$�J�㑶݆�Pq��9�����rRA<g�R|CG���UEi�em�S`
mc�����oT�e9���x�����SԎ�����#��������nW�>\;=�*X/moS����h� ���MV,7��Pk.�¶�������g���5��W����f![�F�S��Pv���s�T�;��xI6� ���a�~�&����#��S:SK1�Y~�6w�Ha�X��T�8\I��I��6�����	�0�2(��߁���tn���ܼ!��,���ߢ�m��s��O	$}�bo�$��^�� ��˓�I��7e�঳�����P��n8�՗��]�_�G0M� �/���oҨ/��'Sv��5�llS
_��)�=�a�`��M`��hCsvMV�?�[���z�=n��a��Q�е'4�2<>o}�Zq��VC�,mq�t�X�*'z,~�X�?� �5��!�����e@)+K�V��#������5e�#2:"4%�C{6�w��
��jX���VL�v�7d���I)���F��pMTy�#�sNpd,�������O=�Q0��'��Y���*!����r�Xnm����C+v��*�b��rc�.=�Pp 9wS��(� �AԱ�r��"�b�s/���t�?�l��j��Q>�����s7'(߿�^�^P�S�M�����;�B/�0�w1�o���V(&״l�bJ4!�7-D��*`î|2�@�Q�J��ᏘH�S�~*X)}!�?~�m�Lށ�)��a��я|�:U��x���Q����g6'3���#���\�M!]��G�v*V����G�l���1��ӱC;�RЊ:�y8����W:q�G�ѯ��Vޫ��D�/���Ei��;�X����!��{j�U��Q;��� X�\�J�?�x���@��؎�]M���T&u����a�i�(�oWԯhοں�~�#�t�����{D�jm ���pk.��//�v�N㾠�~�e���:���y��]mdN�p�Sa�z�~��H����S^(<v��<� ��L��c�#����4OBB��w	$;� j���W&�3[����}���m�U�|�S����(���"gI��@λ@׀c�G	G��x@�.���/��ͺ#u��N<l���uJbnHc�]�߰&<�Pכ� Z@%���{����`��Ԙ]/rgjFh&��т��$W�ۏ�<�K�e�/�{"�d�z���dNs+���{g�֜��,%s�$�e*\�V�F�=K ql�.�̃�3�}�R|��F�!8P7�?Z��{��W�ц��LRQ��>�`�t�x������vKA�������ce|��bO��L����������Q��38���V�s�~�V��H!����p|��
`7�ұ�@��(���&_�}|�;�$P���t�D\�{���j���4=a�ᯎ�,���}�Q�yD� p5˕�?4r"! ����WDMf�^j&ĉ"�4ب ��*��D�^����S��+ߣ]���ȉ

r�,�L�ڤ���ϓ�N�l���]n�	X��Gm������C���V���gI�j�Th�6��e
f��;+J�3H#+*tJ5bШM-u00�n<��m.�A�o�]�zMtK�M_u����
��~}�^��77L���,)O0v���<N����i5F�-y�~����1\� ��j�&8e!�H<�y��3�i�e�N	�[�դzl���?*�޾o@�a��;(xo#�6��K^!#]�R�ַb���?�D�O*C�.b��7K�]]}�&���EZ�f&4ӹ���/cn�����fBE5fn��5 i�zʌ�C�5�w�WP|���4����[Î�p��պ@�V9~[�PT�xo*��*�Y��@�.�Br�۶P̎�K��М�j�l���p�j��P�kw?Y�k����9�Ī'�0r\�x@LK2�~�хP�;QM�N�]�݃�?���k`���4ܳP|t���mH�K�VvU�U2��?A�}s*�pI��|�-�c�{:涽�B�|0�+Ǣ�E�<�ؒ��Y�� ս��(����!��{�\�bs�Ͷ^�ځt��I��M^��>zJ�ۣ33�9�3����`$'�ڶ��n㠰�W�VE��ocW%1	�+Ψ����� F�0��ڤ63Z�^�ck�D��ےEЬ�-����G�|cu/W� ��ԝ=���f����g��������Ȟ�W�#����D�c�����H}��;�ҝ�G����:���-v��))�	��.���ZC�߬�h������h���C�)�?��Qu�wPZ���)������ʵ����JT��Nэ�A�*1��1�ƚ5�7�4��'k:�D�(�w���qP�����\�u2�`����44oJ�>�
I}�yRԯ,��v����T>�U��q-�+��2�R&
���8a��;�>_��a�M��3OC�����=���;�h�Wl6\�gJb��2�znY��l~=A}��BN���[���P�~��I�]��Vf���O���Szb�D:%hm�zE��o;�=Y��*6l���ǂ�b칉��Y9�4�3A����I��� �P�[�2�"ʷB/ǯ�+־�b�6j7�q����A4u��:�"z��ݶ��5@d�uۖy�}��xY\���~�`<t�R]�U����Z��xn��E���Ax���f�įyD�k��o�C-w�ň��?�9=;�9l�U�(��
�������$�	�ɜ�|NIU
�W�l�D���ŭ���ˋ�p�3��cx����S5�K�\�'��o8�ʥ��^O:��ߓ@#�������&�y]	.����j'?�[�k&��▨�J�O1��~)s��b�F��H�+PH���AFw��C�2j=҈�i�:T<7��m�I`��J���K�C�؃g�(��[��g���7$�)8׳��T9/��0�/&>6�j��29��&۽�i���������;ܛv6;��ܴYf�.K,���=�Z�.#���t����&H�^�@�\��A�zN��_���:�1}f�ÈB��C�F�_ ��.����"1-�iGӺ���/h�O����([��q�V���=��>&/�P�tI�~Ʋ�%������.hY���l
='����������y� �Q�x!菣T$�A����9J��~<qO���`]�M.�jTp����R.�1HS�S�ho/jL;�z��"c���Ԩ͝�"��1�$Nє$�f�9����`�R"�vG�Q,�����=���gPf���x��abNL{����m)�)`hx��(���0�δ�7K����s+:oY�T��j'����$n[�z0��rD�M���һ��8��;���Uwn%��s�wCj���1�*����6x�C�}d��/ȸbF��&��#��/��e���u�o���"��a7��X�E����
�a���w?(��1��� F�]MdT/r/o6�\��tn������P�0
I���ҷ ��=�8?��.� �h�8N�{N�g0x�aw�lݗ��8R��"l����#��8��l�8��:qb�$3��u�@�P��p�BIP�<׏@1�K���1*wM�#�
��Y?T��b�J��	7����D:�Vl�\6�YZ���e0ķ��x��Y�<�<�b�5�vc�y�����!�uY��)��W�e���8
Y�X����	�'J��et8ua
$,��=.�q�8YK=��ꒊ�R&WҞ�����ϧѵsO�}�Tj�	����w��]��@��ei���-��@hM;3�֞�-ˠ�s{ڡp����r4���׮.�Rcm/�����u����X\B>H���c	��	��($׆,C�@:��Ɂ�	���*<
,�E��5����Q��<T�߆��⃍���/'Z�V}L\�Aj�RZd�9�J�� �_PФB�����؍���+�+���@()$TH�#��"w����aW\�6�HSa��c���e��΀�T��х6}���#i�1�i8���-
99�����PW7�9�m�0�J�����vB𣭤-3,u>�_�c�N�uL	��i�B����Q�s�Ş�'���MF��I)Y��:D��oL�O�kr�-���u���ԓ�}~*���A�)$}9�b<BI���)�o��H/��Am^p��0��@�p���0>4�L=t��vA䔀���5�~5��Ӹ]��i�gS�e� x�i:i��-��l��Ρ�VW@xrI�п�zʧ�vCTΒ#d�KepN�6=�!�܄�����;~��>,G��d�O��rDhY>#F�d�zaOݫ��j�cC}��h^�q�'Ԫ���:mW�c1?l��G�w�;�(;��}�����C�_L��y�L����
�~�Yw��<L�ph�Eư�c��,c����@�4z�֌������Cb̿�e�����0��H�m�����[m+ÈΝ�j�\����6�E͘Z�ϼ�����L�fs�.�vf��� J����ğ���x#�ό"'�\p{�����s	��K��4+]u��kB���ֹ�?�k��-���K�[��q
�5P˻�Q]����$k}7;Xd�M�z����F�Qu�ɔEb������S*fHr�!�\��
k��L=��R�qV�b3?�mjN��{Tӣ�*:͔R��5��^8��xT�]'s+���pEQ��0�4���8܍ѵr�^��3lK!��o)�G\ޯO�����#w�\V�e�Q?���=q K�b���%`�2u�㪬Q_�E��AJ����r�l�~��B�+�y��m���=Mp�@y���sJ�tC}�x��vNn�={��-������`PW@�/��.y�>��J���)Qz�����y�Z):�~b��"��Qʦؒ��lS�.�Ty):���3n ���B�usO����Q`��W�0_�_�A�V3E�;�~�P�E2Bj�Q�ŭx���Lk���x7�4���U�������
o��9�"y[Xq�H�Ht��C���'RpF8ت���e���O3�=�sU<�,g�sͻ�Ug�=�;=ʤa�JbD����Hf���Zku�g��s+	V2�����5t�'@�2r'GgEw���D�p�0T8�v�L�C]�ٰc�*y���������8���0�8U��v3T64�L�B�>��C&Wdl�%Fޚ(�^Ͻ����	xz(�<H�!��~i-���w=�����8N�GD��ݛ=E��o��C7�̽�mFlu+RYQj+{V��������6K7�y�c�l�I)�|�FC�^�4+��K$L6��Ģ��p9�܉�W-����{%�'����OȂ]�1R���,GU�K+D�U7����<̽NP�6�1{��+L�Ts�x6P����S%c���bI�����X�9��:�m�<ѡ��8�'&�u���=��wK�r4q#��5�N����`+�$-I+�37�e��~������b,)5/��e���^M���3�yD]ڽ���;ޖ>�8HLD�!T�{��,� I�Z��:�M�`�����U�c�����d�*�1>�{\��G���ɬz��f�gH�
�����v�_/0��z��̓��,)���UG��"X�>��	2�i-��9����5Ɨ� (���@��E*�8:J ���)�)ۖ<έ�1�n�hgط�3��&/����|�[X����HuzL8��.��Q����k=��&Y��;��9	��_��kϢQ��l����*��%Wt�i��T�%x�z����@t�k�"vmo)ʕEV�%	@�jФ�z=�L��{W��vd�h��ٜ&���LH1'<�S��akq) �5(_���[4,�%��9!vT�+��NU��8�:�?/��_�W���tj���b�����v�{�=yJ��qkX��G�^��a&�&��բz�κJ�s�_�e@���uW
=� �r�q�I��@|�ty�MА�ɣ
�!�j93�{�K|���
��8��vDR!y���l"I(꓎�1m�f&wP�=�1�U��pN�(R�*{���0D�2pd�\ٱz�����Ҷ��	?�ӂ�IU DB����bi�W'��-�si����f� #& A$,��7*_6��6��{��װ���E�/�����7	��3S�J�׹��N�H�3��0�wMX�%o6%����<��]���o�o��*��Y ފJ�>���0_,�Rw��oI���\�s�M&5��cմ�ֿ���b8w2$��]�~p��h���{N�w�?,��-��{���&���~j�o_^��@έN*�9�����w�����ܦ�h9���4��	��1��tx藞~U蘌]x?%-�f�����ѝ���\͗����ꑛ��>�0��ۣ�������*��� ��W��A>�vX�:b�	H<�2�ŝ�>�8t�d������It������)���S<��`��J��vldC�������-��	3��$X
��2@�pU�q��ʂ
��W�N*�3	�����oĩ8ZҼ�¿�;NjvC�����`�l8��e&O�H*B����>�+s�L�w����|4R�uʰ�j����s,���$�L�.�mB�n�r��iR	g�L3xӇd�	�)L5��2�+���bk���@�����Nr�?a0p"�g��c�W"�����D���l��ßо0�-(�������0g��:�q$=�P��AS��N��&	���Fh�(2g�k��ǂw����ν��T�%[��[N֪�������iΟ.�3��e�P���7��i��[*�����f�F�V;��"yk�y&m�3i�8&R��X����ᕯ5W~�TV���=)M/`�78Ix������j�Kէ.D9�,����P�)���QJ��D>h��}�h��s��'��b{�T�3�ީ�'��"p���X��Ĕ3D�~v���N�g�T.R���E��L��c#�ه9_/y��ׯv�k�`."M�LY�i�i��u���kj�7����dh* _��S~W�.�0�:��Y%���O�Z�ӛ��{��pO7N�/���H(�i�%K�lO��F�������V����{OA�!�c䠊R�l����~"�����v%0�zw>�a�@*9�i�Xt�
�6H���5�L��J'�kJ�ۼ��!uz��/�vc�������f��ٽ�J����z�Wg�'7!f��r�7�f�k0��p�������x��`��@:�TA3��	u'Ө?�;�.��QXd]��Q�K^���^N���<��f�,� �Z"('��AO��ak��v����_~J*>S�`"�1!�KV遻��~�>D�Qs��	�ҋ�ZAAP�,-E>Ż`�i(y������K釸�BDG�'gG��\�[�"�bt��DX�܋K�/r«p���F��aK��-2	���Ʊ�^�B�d�z����a��_�j;1�|�Ԁ����jVk�^��p@�ĩ�d/���l�I�3��A@��2r��h�'q���*bܓ|_=�3K�������$���<7yR"2@3@�⒴����"��b��r�"0��W��$x�����Z�q8�m�K;F��e�����O�ILe�ځf�B
R����B=�Yq%/�)Q���0s��"��%P� ��_�Q�fj̓�ŉ��>���!���<r�a�c`a�W.��X3�u�sh!���^8̷��R*��-YJx�G�3�mй_��g,�C Vj!��6���ԒJ���aeB�m{l�/���җ\�4'��W5��s��<+znԋք���N;ҺXh������8�Yx��fZg����iY3j�Os��t�F-��������V
�p��ؾ�)���$E ���+� 
k׫���t3����ä�-�a�A�m��:�}2@
_�o�n(����X~L+�x����ޫ��H��3b �Kk��p��f����1JqЃ�{��r��*	�#$��7�pu�G���5�G	-�W�8�8t%���G�8#j�ս@�ԅe�V�O��P���p��7�Q�V�D:�e�@A�;��`�=�j�CML�0c!JǏ@^��*Gd��v�p�_%�~�tN�����2oG/S��"wοDF!<��M �soH=�q`�;I�c���f�d���I�nt������N�8&�]}�v��=��v��J�9Oɓ}��XBX�Z�[�p�mz_	��fk��T)�J;Vaz�ݼ�7Z���t
Xx�B:�c���|�F���l%����$[H��0��ީe���6�|gt��%�RU���G����_k"��u� �u�):�����~c�j��(��co���R�z���ʠMB���f���P���>�U�MO+�n�{�{�֣�s�9��k~���5mۇ�q�1o܆�7��#��핵��q�a�RF�����7%`e���������dv��ڊ$���%������0���*��K�@{��%���1�Q�AP��<�[�$ e��A�Dh��nߙ�$_�������IHs��ZVu֍ �f�oG��دW	����ߙ�W����]��A�8�!� �2&�F�5�'�?�y��Y�z��vdｑ�����:_�aGj���W����ۘ��!,�y�ysRm�DXռ�{��soœ~rP��'Nʓ^��+�;���Km���)���0N^����t�y�񍅋�D���'�h�q�K�ӭ���?����'�l>l���1`�<�ߦ������X�S=f�*;��q0���N/�`Jd��
��W��+[��݌B@�m���St������,E��32-�2gh�\d�h� E";�/XBSb�'���m���c`�1��N���sK���aW ������ě���t������b�Q��˨'Qp�4��V�B�י����T��w�̀?�:�)X қ�A|ZL��4Ҷ�'�x�#q>5�Ji�F[�eT�B_!:�ʤ5j�EJ�Eς����c��� 4J[n��Z�j���e6.�B����Ї���-��c����X$`��@��[�~���z�oj���mZ�eNC󣽀�`�J��_�!Z����μNҁ�����0��(VfZȧ������v��Y&{ۭuYlcwD�|Krq���Q�r�B�ݤ�h�!�3�6���*G�|���fyiε���}�gT��[���F9<O��U�N_�Jr���wo�V��n>L�Y�a֮��:��� �"DH���jw��d���q��("r�ɞ��L��+fզ�Z}=KN�rg�Ra�v�;G뗠��9c��Vk����KN�Q�s)�,����&̑��r.j	$\����_��36z9��ƴ��|�����)v3���bf�zQ��* �/��x�1�@,z�g�X��N:���}.�����Z|��;�ݡD�%�1�:�K��(�O�0N2?�/�{�xR~\�<�tL�	����t��$K�,"��8��Rτ�9�� ��J��ə2�<�q�\�%��x]l���rK�hP	;9=`�l��2�.O=WTl�Λ�"����1�ҫ�O���S�Ohm^�g���.ލ����ܬ����=��!(-j�}�D>�(��K]j?l Wk�8-I�a9��Ud/|�.����u)6����q�8?W?QbQ%!?	V)XL�-�wC�W��5i�u6��LS�`O_�C�^^����Z �I 1jѾc����e5N�?u1y�c���0z푏3���n�����]�,ʵ�wq�?_D{��K�E�j���b�q^�/�J�o�1��~�T䎍�'����:�������Η�T�� �<�Էhm��J��t,��b��V�Gp�8p�Q�$���¾�n���Gp~��I�����RCU��z�^����Q
�'�A6s1���^�4���u�U �e@/��v��E{hEw�"9�l�\7(<���,R}�5��}*�o�S����9H��M}�໨˺�c���v/}v�ծxO]ր:�pK�#����vo[��e�zO���ؘ�	6��6L�G��$��Umx��HG� ��6�����i����;a/�����J]��	e}�D8sY��W��vb��6pF:r�1ֶ�*(�ܪDgz1�G���d�i�|�Q��9BguIb�y�Y�wY�7���ԟ���L���2�`!�V�s�$�lY Ap��h��ݩ)��׫E��I�Bs�9�B0�g��������s����m�YUH�.tG��:h?Ά:q��MQ.a�����/�f�����{�b6YG�����6��d�ֺAR�M�m��i��o�Q�dFwX/�18�~Ce(��xVB��D>oC옼�R����\��Zsf:��Hp��K95EPךځ6��S<�%.]ȭ(�l�Щ�&Z-��#�W6T=:܂Aq,�l�{���\�󢉶�@���T��-9��셣��?��P�Y�|��k!�Y�F���l1a���}�
]�9\�N�~���&F��8f"���N�Ǡ��Ԏ:�(|�u����D��[��ڗq��~���)#~8G�\H�����
���ȂU���B�Q	-ͨ�
�U��ÿ^3�ѩ�m"t(-�)F�q�W�v�$��c$ _���+H���=�5��waC�'�g1g�.�ʑ躿I/M܀F\�>϶��t���'M>��_O�����I_xw����{���_�ʱ�0�_x��&���8x�ň�	8�o�C1}���]��3��ꢣ�1�%�
����#��	Y���R�!t+��$�`�����&��XY�� N�'d�$�h��[��{�18����`<�������-�oq��?K,��=e����ѻCBBf���?�/�x�_����"���	E�U_ޡZ:�UPGZ�F�%8�M#�5x;���5f=�<M���bg��m��j 35y���nc
gu�əP�o�ƣ&�K����ޞ'��wr��g ��9Y�i0����+2���"m�O�Ɔ��ЉR�Tkl�H�S���A=��4ch[�1*�����=U
�'ڭn��%$΄z�ōw���8��+ׄ����� 5��{s��G$�I;֔�wZ�T󇷹(?�?��䐥t�̅=�B�O�5Kil{J�}�4����;�	i�`��0�s'm��)U�=��OQE���/�G�r�CL�ӀMO?�� zĹ�ɂ����0�g�lT�J���0�ad�(�`�5�Jk-W�x��Wm����e�{���GW�gɛ�@�I�kP[�w`R1�=M�۰z��Z�-��r��3��1�{J&�� ;���%Tv�<� ՆuN�o��sh����^j�����߂�r˿���u������}���p��#L��s�7AK<��5$eFǡe�d��,W���`Z`
��+&(���T*�z�Zc�͋���ﰁ��3��-q�G)���%PO�>�4����6Q�o>���`�"`�/T�e���l��iZ��U�KY���*i_�;(�i/�x�Ӻ�b����a�譜�s`[ݲ&�}�S���<�-A1|��3���]��~�o&��po�p�t�r�V��Q��? *��r{:!-�%,+gS�lo��[�S�w$��"XibQ����'���0�e.��L�@l�VB�x���?2����h�C�Ě<�ėJy>��#79����+">��m���68�{�,�+Ţ���^�#o�Wߞ=Ělu�~P����N&.� ���6.|���2���	��#�(	S��g�W�g����4Q�]�貖�����\�)�
N`c�G���b%>��w4���%iV>��v~��{2A����Λ�5l�����	>��^쭁+�_}<�����*I�C¸^�����9��:��!�G�_ȧ����3nM"���1t�"�	0��(���������3��.�U�H������,���B4�q�2�=�!��<��6]ّ] �W��M$�|������������伔�f�����⌉`{3�̕�v��/;�,�HڒY������N�h��il�����vK���%���B��d����M�����A�����S_?2����*�N!D��}���¨�~||�}~�͢M����S���$�m'Ų�o��s�|�5@M,�O(����U͸��4|����U�O�}gi}�=��6Q3:��5`�x"!'����Ԉh�!��kȇ\i���1@b��/����OV.�3g�d��ڥ���8.��n��!B��Π�
����o�bIhov�.Mz����^�n�^��ڸx�C�z��H�E�~�>9c����cgd\:k����r<�4%R�M��ca��#�	H��$��Dȍ�S���!��D����j�矤K;2,�7��n,�f*
v|/(�6�рVT,�PI��ؗ|m+�~۶ﮛ��/S����2��B9�ٶ̊�Hx�c?}d �R�jQ�$�C�ҧny/`��_8b�ߣ
�i�Unf�2￱kdW[RyM�t���O���v�ҟ�]8K)r���Hg8��`��}����u���z��`!%8�TD�u�7C.�v��C�jb���I=eպīܮ����>=ԧwq[����4,LFƼ4������s�:w�Ƕnp���@�l/AՏ:�7�]� ��ZX�hU��Ӥ|6��Ѩ2��DR���0 5V Sű�p<T�ǩ��H_9�[��FLD/ˮ�Ed�3<�J!X]>1/%{K0���Ѵ� 9��	��CܭF.Eٮ4�ё��^��̎M@6J$���lK�#�!&=?��H���w?�d������PKx������~N�#fv�ط�����&�Q;h۳#��K��m����ԶH����h��n��g�0���bT���!a]3�� k�,=;��#�`����f
�eN�#�!:Ox��zيS8�q���K?,�"�ͫvw�s���߂�Z&;��V?!�,� '�^Iv��Q�l�Xbep��Oס�\kn�+�լq�o/J1-W�䮌W~}�y�,kWQ��.UNWu��8@�ЍbE��s�v�'�E�����^���L�|=�A��]��lsʯ����+�h����80�w���d�4���}����3�޹$4���<��ċ�
�͐J�%����ƃ�E�_�/��"`ru/w��7ZZ����K�Us���Z��T����Km��h:-%M� �)�$����ݼ�8?�D�&+��m$Ē���� (� S��Q��S�-r��)_Bu��Ѱ�0Z�0�Q26}~֬RBi��j��4)�D�(E�r��#B��<�)f���+wG6I�㛊@��|� �^���ՊkZ�>X#!޵c��z�5�����邥�r���/F��[����ׂ	����UÊ b�������op��}��X�~X�`F�`H6a���K�0��.h.6�����W��&���5'�t�/���ۖ�.��YjP��$g#����Bݔ!
(�����Z�n;�����pVC���[b����S�z)
9!�P�p
Qf,Tn?��gJt��40��>��H.b���w�a�S�&����K Cۇ���k��v�� g��A{�x��u�T�g�M��Z�I�f����lR�G�>���=� ����c���0 oS�QK�MVQ�����!#N�����^W� s���2���W\��?[���P��o@�bX�2�K�\�I^?�QRw�]7�s�ۅ��4������5�ؚ��Ҽ�(��*a�W	�D��"ք�H� �0�kݯ�C�/~�J([9����R�&b�g3,��V�AU��*H�tb�=.b�����+PO��"�f&c5Ft���m��������/s�~�n��ه�U��L�4��k�T�׉�ނ?+�S�����Ed��&�}�y���Ðv]m�=hJ�� p\%�2L��L'����(�!�V�<Wz+g9Z��o�̂f�8}�|����
1��p��^���(�V���A�L�}M�J��BaJ�4ҽ@Ӿ����I�|R#��������#�.ٰ(e`ʗ���!/��?�!�H*�Wf_�fl����ݦl!��}�_�_�OQ�S�%X*�3cTX:-V�_uZ��HxCo&I��D!-�'�(7~�#�S�d^K��#���^�����2$�TQa�:�0^�AQ	�[ǩsA�,�U6�Z�4��iU׊���g|u��WH{`��;jv_��c��u���sy� ��[0V��Rs,j_�Sm�z�����|m��␆�U\OgM9�A��%c-!~`��aHn�D����%�3e.��z���h+�����(�~��L�eI�8� �����'i�kR�V/�Y��x
���PU������?6-b�Y�w|K 7E�Rg`�Iؼ��ݙI5E��>���� ����w��:'"Vb��sF��>���i��1��0���[`�!�q�"�R��N�wqd���-��O#�MCS��k?��P�ͭ3�u�@xئ�o���o<Fl.�@|��*Qmr��ż���@B�F]f�]��-q6��B�k�<CH�鿡a{�и��;M-'l��.+.i4N�mսU.�����V�C��\�v&�U��"$?A�x�� ������ Ai;FW����L�ޕ�W�'`�a�B�L���3p�ER݌�c��y�
BZ��a�Ro� Sz�oQ��=N��;	Viw��v�u꬇GKN(��vT����g�t�`m<��e��S���
���8��%�<ݑz��a�ɂ�=���;9�!��V��3#1��kA��}�#x~�XNH]�z��%,8��<��Kewܻ���UU�M$����=���Q�E�:�ﺢMjÔ�;-o�S${;���5-u�a�*�`a�n���B�P�G�+�6vI�#y�����n�p�rc��d� c)qT!��j�Ǭ�+���2���'J��o�@���}1�!v��Ͼ��M��7ѹ<�)����j'o�C�
�L�4�;no��Bi;��5
���U�8y�^��6�~|TY�M�g�0d�C���U�@ȦL��Px�d7,�m�uz���*"J�ߋ��$�e��J"�����`Ќ�I�Ek��[%Ã�xX�HrMdT"&Q���1�f.Sڝ:�|��SUH~���o�Xr�l�v�c��sțn����K�ȡ�E!^bkf����_�A����m���}�8���ٝ>c�mw��w��J/��.���x�BWן��S����u ��>ȗu�-X9�On�$�`�����N�-�����
v�?˸d��{�^&z�璋Y�(�[�*u�x�6jRy�AK��H��kbz8��g-�B$�T�Se�ޚߑ��[)&�!�J�`:m�r��D6<Bu�k7�8p�,��\C���#i�L����֗,�_�`�Y$[���>�x߲��SU�-U�7�C�C�x��Ԟ4�=	�h��.],��\ZȢ�Yg*A��!�!���Z.���׻"&��l�0"t̸���U"��)J�#?�B�gHT7��G[٩�FJ�˵�x�2#y���as��+d#��*��K�v>c�T�A,�w��y��я�maI0T����e��չ&{��߷�oNW7���Ӷ|Qu}O��\����[TO��< �E�O%[���-��kF\�l�Lfq+dG�}�>7H�p�:aSW*����d:����M�z���C����x���ӳ&�%���g���?��r�N���!E&���oJ�٣�r���} ��a_�>R�i����=��eF9S�O� "te�R����DV�S4w�΢�BD/���-���@q�6�,L����+
՜�5qk?.��^���?Ą餆Ƃ�z��)�n����7h���h[:�Ҝ���x�gxfNt���F|�a���a�S�SM��!��;��^�a�JHR����� �	�O�+�G+��Z�{�*j����j���>r��T���Z���"���R�]E�]�c!B�5h�hn`4�
���X��*�T�|B�Op���9�������c�p�Ҕ�]ˎȫ�bafkMa��s�!7h��XU�t��_c�PX��b-Dw�����HҊ>u>���l&�S�׾����p=����뭿x�� �X�Jv�`�١o���������J;B˒9�.����S��5I��]_���p��[�%�\�l�J3���ټU��K������;"��mX}��n����0�fQJu�H���M(|W�>��I�9(	�ăRi-^�_��c\Z�:8߿9�j�����Y��+� C�48ؿ�Ŝ��J�'a�%������^�]v2ygo�~�@�W��iv桠�����~8���Q�f���˦p�c��s
k�LRs�]d%�̒��%�ҏ�'�"k��|@�TEҎ�l�<�Y�0�{@�m��4;����!G?�B]�������ey^
c[�&bH���fA�2��Q�6S�ƪE^h����I1��<}�S�*���f+��0������<=3��۠x��s/�@Aʻ�P-M��9I>�wPRq��/�0�q6���K	���̸�w�-1���w[�S�
�HO�z\��xT���^���b�G�ZV�^B�,����҅p�t�~��D6:���
^x�W�Q<��=�ȅP�m��9��	�7	�f�_X�ry�(),�K�b۔��6�� r����9�/6H�A
��lUT��xX\ a�P$gOI�O����T�$����o�="��y_
3o�!K�Ք`<�r�gw�:��jt1��[�+��ƽ����a���=��S�|%ҭP����s��j��/�4 ]���EO)������k�d�Y#U���2!*Hg�(��uX���H�b<�sȯW�x�}��
s�_<ZD�� ��%%	A(b_��5��|����}� �;+����ٺo>2���c�I�x͙2JcR,"�H��LMݾ$���s�i�\f�'zǮ���{�%���.�����^�V���[��S��
l�ŉtɞ$~Z��	{���nҙD���
�������J�[���x9�t�+�q��c���NV �����xل@JV��'K���N�4��J���g)S�U|�b�>X��C)�_�UJ�1�D}`Ю�B���| kf�́� â/h����T[�y�2"��{���F9j�!w�d�E,Cd�î��,`����Ω^T���C1@��A������Y��}��7�]P/�WYZ(M�������n[\�s��t3 ��F)�3��>{~�z?�>����+���4�V�i���g6z� ?e��K�z�Q��%�I�?�ߓ�o������ӈ�ޭ݌�h����ᇺ�s]��@!��|�GP�1��X�7F�=� ��\�q'�c~�o5�WBP�n�|\�?�u	d�O���)*0�Ir�2����ֶe	,I�I�V�Q��*�� �TsW�@}�vH�+��q��ە��Q'3���h{w��]��̻��Zp����wBj�õثo�D@��=7T��j3�o�ZI[.3�pI2հ��'4�r�5Jb��5WC����	�F���6��݃�d?~Sv/Pl���LB��~�B��Z�����]��\����ҕ)԰�n^I`We	[��=���"ԏ�K�����cI�m�MeđS]G���>�|	�qb�@.��x'O�\�'�.okR��h�t;a���
�Y(jlA��o��37Q�㤸ũR!ƨI�/�JJ]��ڡMbw_�~zɮ��|#)p��<�rT"�4�4��J?)#�� �H��É�`fR�7�B0��Gw��6�z᳟)*AH��1R����G���~�6.ǌ���պ ��Ź��!+L�Lc������ؓ��V�`e��6�jb��� ʝƯ�u~F�)���
vKHM-b��-LW�p(;Z�:ډ� `�{�MϞ}�O%�1�G�1�`7U��_��і�r���rs��/��J{=z�wU�@a�-�tc�-O�T䳥?]j��	��xV����|�l�����FI~0�(܀�sN ��rI�|��JsN�E�[�W�m�.�)��@��v��N���ĉ�hڃЖJ4�C���jMC�>b��W��]ۘ���y� ލ=�a�F.Qc�}_��	�rW���� _�5�6BB"Sv#���=�it�E�%ߑ��h�➈��:q�t��S��B�S;C�Ϝ*��9����<��9��ל:G��o�^N=y�%�t��I�rU��2_�pm���F���v��AA�������O���A��x�2]�Oȷ~��Ek@�P�D¸{i��{u�������!rg���EDz�\�h�d��c��������~n��-K�\��N߬E� ��[$�*悁a�?�񨟨m�X2����aO2��"�B�saxh����� ��C��؆�k?v:ӛ�|"A�3}��!��V=y�m��b�ܫ [�=&�̒!&���m����,��1�?�i4Q�3+oKeW�+�'�Tl�9��[l_�T(ڏ�q�tpGi��͋�_p�zo���PU�4`q������錕wxED��1F�2��5]�r7�*3�����[;`A�U��3p�z�z�!��s4`,���[yڶ�su�	�+�ړ !_'�#ę���U���N��������|)l�Y>L�oҞ�"ui6��I`?���2��d��a�+� ��i��`9�OQ(���N��&KkYw$���L�~t9���;���b9lߛ�yj�e���H@��>��~�h6�W�*�����Ԙ��ʆYF���	:Eh��og�ц�2hd�O@�Ņx�� ������Mᇼ������Y��������f���[R�޺@����f���.�(0��м[�g�i=����V���P\Bq�Ji��} -�is�8g����=�䛜ء��P�6�+<3A��R{�Uݧ��M��SY������f�@ǙpƝ�2��/��&�~_R~�2ADғ:���t���܈ǭF��k|$xj�o��p�����R��yln�-h���b~�,
������QVb�j
��=���j�Q{�J������\����!���\�����S��nN됟,g/��,jz��
�K*n�������H���y
E�>r<.A5{&��;,�{ .!U!���߲#y&�E�����'n`%����[����*ϸ\���ڎF�#1�M���"���1F.${W�󶌩n�L���d���A�.��
� o���	��
��=?��lgUn���Wc��K#��)� �2�R���7�;�� ��$�fr=�rL��"L��7���!��"91X�~�c�e�w�ё�;�8�K�Q���γ�.AF�y�ǒ|���zH��=�*-Ď�0����� �F���E�������������8m�ͺ+<�P�Jz�%�ƹ�`�n��Ř�T���~|&W%mIH�)�8i����;�:����k�Ϩ����=`<=_��_~� XB<4���O�+�:	w���;?^mm�F�NB�>��p�~�������XP��;6O� ���v�s�^�%�j �0ѩh��C�z�Ѥ�ֵꌳ[_~4��(O�,yN��2!����i���}2^B��n��h�H��$"ͫZ�:}� ޵�]�8'��J�T��tQC��:�����S����]�Z.o`�w,�i�E߁bYM~=�K�w���X�$�c{�ǥ�A��c?��8{I��B���K
_=@ :`������T�H�w1?�kӧ.�W��o3r7�U�a��/����?���A�Z����IiF�GI
p�D#uM�r�_�Ȝs�A#O���:8��:l;�w��|�#V�Y�?��8�׊<c�<�ɦ=ʨ	d�,��ݪ���;n���F+� �\��rcR�bm��Ռ+��N#�߶�`�C�h�h�$7�R;��o�v���({K	f/i�A���{|�K�3AtR��Y��Z�{�<{�]�������tx���|"ܒra,3]3�N���_�9���s��!�<~`�G�b�#^�Jc�>��-���^�e�֨���A)��in�Јs��AwXA>��2z����̐�U;�a����O,h`��@� �j�إ|4*���w�%��s��9�N��4Lx�D@�X�_m����Sg���3��i�ҕ�ƙb;Hs���N0\�#�Y�
L�ˈ,\�%? $���^ӣ0l�
4{:�` ���S��k���� u�Ai�A3���,؏��[>���Lh6�'��	9�2{R�:���rz�)�ȥyr�
���RÃ�=t^�m>�S�'�4�����8�W�Zuh��%I� ��[����5�&,�<�Z���U~�0*�t��f�I�<��r'���8�CDe�F�ӽ ٺR�s(�7���%),�����]������F<C��g�K���MS1�
{w���9�y�]{a5y�k��w�Pл���.����m��k D�	��@��S���#���Ƞ[����%��k��1�ڬ�qs��`:?����f�_�Q�do��N��
��nI���!*ق�c���TC�a��3��=_>�7���mZ`�>g\x�����[-L*�>�`3���
�!'� ���kF1֠s�`�G�4CLy\X��	��|1~�Bnh���P8�e�P[%Ԫ���L(ei�eZ���,�M�bX��7+O���`ʀ�-�:��.5=�'�*�Ei���(�Y(%g�u�}T�#�o 1��0��6���.,v��PX'븗�����mD��X���1����.4�^�y����n��&�Ͷ���O�(P�Z��3���� �<��֪>F؈W|B�e?�������� ��^�٬�,�"� ��jd��r�Qo�1����e��~񪙺�ʕ�b�˰�_;_D���^�ǈ��۫��i�Dz����r0$�ݡ;{�Lj�U��u�cSUVBo/Ңb�E�c[�xL:�������.����z��"��3uj!/U9�������`Č���A~����.�xY���3�餺JL���z�q.�l��(�k�/ŀ��
�W�#p_�9@9�ug[K�'?LA)v��M'�c~��H�V[�F���$K���[��)��^���S�N?���ҟ|9L�&3�ٹ*p����UB�s<��{�1�-�"U/�}cGz�y��(hf�]$��?����E9`�E��K���i݆�+��b�;r��PM)^� ]��H�7��������]�%U�uH=\N2�yr��m�OىG˪��@�^rf�'��O��)J�|�@p>Ǻ�C��.ĩ};F��������	1,��)�n��م�8+I�I[�H
g�
&�0UP�D�
���ӊ.�b��!���5H�(�v��-5@��6���q	"4wX7+��7*�p fl� ��E��/��%�=u�;���܀r��!ۨ9�(a��?��U<�$@�X�n��Q����uf���y�Ɏy����n�+2p|`�S��ύ&�Z�p	�Ojed˗����Y=���ڱ[쀕tDG�u8��$]MkW��� �ZXӨ1���\��K�T�rCC5��c�|�𵻑��ڦ� �ʨ�) ��%Ld�N||��a�w-�������.�T��w35x֨0��Cet������f�W��ׯL� y�?�B{@�g�0��c�f��O]j�����p�g�<ࠎ�S���4c?�=�L�UP��$��~����Ӻ���B���5�^��Z��HL0���j|� ~_��X�AI� ���Z���`�e�6zL�����%��Y������JF�������p�g�W�+��ϣ���L�r��k^�A��۰����ճ?��Ujx��"�DJ�&��d�X{��,�@�߉_�4��Q��g!��,�:fjV՗���7;(D�ٙ@d�mJ��{s��1��e�(�'Dk���{���1�2~P��l���;a&���Ւ���fU���?����Q3֗ȢzV�<S�J^�"_�^��r�VWJT!��E�Z�t��4���QkBW<��.��|�HgR1)���c�
;��9�T���c��;�ݴ�]y����������'���Ui�m����L�T�0&q���/-Mi��M����ԯ��8���C)���C��u
~��ڳ�1������EEH%�/��iK��I�v�Հ���e5�	%�b���'w`�rr���W��`H�dzR����(6�4�f������bAX���p(�ND�%Ɔ{����ɨ5,����� �&6m�i޾��9�3~�j�@�#����:�E���$�����Tp ��4Ż*�Y����5�i�mk(;'��?}5���Q�O�Ds{�5>�Mx	{E�10��^�Nv�<��~�h~$��k�l� 0D@X��݋{��s@��y8r8?<7����dY�	{���1b�+�$�;������75���@?
|��O�SmB�ȌAe;�K`�l�u|���E(P�{<S��0��v1�y#ym�S� �zP_I��f�/������s��c���m@W׮�}�]U�[�D��{/�'s_�����EY'M�WT�W�b�n��>��0����=$aq���o1R��]�	��R��QL҃����i��tx�x�f�,R0�qw���������K�V��dt�r�&��?x���#�m�&��$Ƌ��z�����)[M�>�����2c�g���҅˃�!�*�B�z�X+W���8�$��g�֝�c�QR���*pM-GOY�����͌oh���\j~�p��!!\��1�t���Cm�A�2��F9S�3fD���_X�^S��h��8��W�NQ�8�JQ$�8y(�Lgٵ��m5��\�k]�-�i@T����W��h�}߈�����N첾K$������2adG><�����h�?M��J5���(�%~B��Q\�H�
�ԧ�J5'MS�����a�ע�K	�[W�m�so��P}n��wT8�Sp<��I��na�EA�������d��N�̖P]��z��&�CX:'pG�{C�C�S$j�I�Ŷ1�v��
|�j*���v����k��R����|I^Y3���E�)��O\	{�t�};
���vz�����}�w6������	Z�T�z���S߷&���h'�����?h!����U�,B�(����gFf����/���V>Ac�%�饰&�����a��ښ�~c�9МO!��Ⱦ.�A���b�z@�c�w��(��A���>C���җ��^m=�[��%\��{�h��X�*�t ����X\�c���Lk#��At�c[L�{��	j�G׎�H�#����v>(	,+4+�ֹ�����9��i�~P{��߀�_���}�X���8�� 6/���H�j ��W��E����!��k4��j:h:�ĀK���T�6�v
C�zL�8��(�}TbT�宍�&��C B���}��_c�tC��O̼��s�v���0X�q:�c8��?>���̜j0��S�/��2 翦F�v��mrMH��1��C|2�e�O?1�r��(��Z;0�b�&�Xf���:;��*�z(]g�)A^���obR;
_HN��S�1�t�^Dd�UΣ�t2�NYabKܷ�],':�3������E��;�����h,`LS��(��%��^�y�rA&�`^F��c��v�)�6�N�ZP	�e��I}JQR�����t�/�hP8�`�5��Oo��
���]+���7���, ^b��3�TD?`�qʄ'|9m�/�E�R(����F�!���f3��o� �4�磭�R� Y���9D��s����7S�Ox�H�_<(���{�BzG�W�����-p�\lDM�� pC�8�����f�󼉐2�?'S�@wR4�θ�CN
o��i(��ܿ�\�����.A����2�[�?c�[:u�d�J<��~����x�B̏����{ZqwW���^B0w�b}˦c"UJ��q2S����GH���G�m�G�2Z���������]&_ǋ3�G�+�y#��e�"�B?D�F<݈Ә����'j���� �Y!��}��&�����QF끽����rK,e��[/�H\�C2Ӹ��L����EUF�=Ǌ��}o��w�Ge}��O��P塚�X ];�F���������x���ISq~F9���7
��Ä"$⑏��e�jC��lQ��(��K���P�i�G3?ೠnK�L���{��I�-���X�6�*�2�9��Kd*��+4$�ne-��D��ek.͌�C)��
���\e_�l.���u��@�(�$9�Va�GÔ��ݏ�U]�I�I�ৡm%�q�z��pҚ���9�P�$k�� ̱�3"��A@�e�C`hm��o�х�.�ٰ?�w�}���4���l���,��o,���L�Ce�1�e����,?p������>�z8mP�d��ǬH��j㋫�d��s�뱭u�?�}M�G�Mx��?�����x�
_�D%��7��&�X?�.���Z�?�_�r�l]�.�����XɀFM��X�������~��!8�T!?5�oKs��A !���F}��`�C0�Rzӟ�C9��Q���~�6E��6{CI�!^S��f�]�;	�����SB0������TB4��TT#�d�;ŉ���?��9���#k�/��C�*v� �&^��O�8��p�e�a�������RD��RnYSR�_um� ���j�G���$���j�H�?�bU��L����?���t*��s?��j�{
B�?P�{�Ǆ?^M7�K��+6��pX����=4���*�6���EY8��2SS���`��|�������+E�X��iw�|K)F�6�.<+c���ҭ�� ��ޣO$�����ى��X�K��ȝ��΅��5���a\HW���u���\��Ϟ߁N��X��s{v��{�g���xǤZ��#�,��x�6�Ҧ�5��԰�R��;�.�Qr��H`R�Sإ@s$���#B��R6��Vj�=Ȝ�cΙ�-H�gj×�L�^܍iM#��r�wq�$%�������j�-%�[�䩱o|��:�_bk��
W�¦ae��i͢��dZYlt��څ&GP�A-�> I�U#1��>�LÉ'B� �����0S�NM�6c�l}T��>��9G�QU0��я�c��5a5	�̝O�nAѦ�o(@��9���Η&�[��#��J?���ȍ6~QB龱C0��?Q���曳>`S�X�3�2ouSa�PxSK/U�$�K��$$��-r9��{�e�Ae0S��1ݭM*֒�mQœ_��[T�_&.�t�K2/�}�ef'=��R�x�cWn�t\��T��MR��j���m�>a�z�+����!��kDlt�����=%�T|w3��ڠ�#V#|ي��ꑔ�'�d3�0wĩ��X���`�r�B��Db���a6[f~P�⒯��א�YBu�YY������J���|�����<ªa���檋E*��-�_?�FiYeF����f�u�$�~t|3���0lܠ�Ai�I��KW�s)��
X�3N����qf�ZY@��a�o&����%?nHz�+�92�_�_r��-P�28�ǵCo�a��>��%����nf�G=ђ�{%������?v��k��ܱ���b�;�7��y��NL�j�1��mx�N�J<��'Nɨ^ڰ l"�SC�0:G܀	�-)������ԟ[-�eN��O��I��ߺ_6��\!X���0]�����Y�vV�Sytp�HZ�����+L��
��V�������|*4���R}��P�c䊧1�8�����]8ܲ�lJ$��-5qv5�k9�=y�F8�0P+�`w�NH��:��us"�#����H_�]�ub�xY�ޮtD�S�qV��j���{JP4�v8ϴ`���ȦLz��;�ï��P��Oc�fk�Κwh��]��-Sd�rJ*��q�㒫ay�f�>����lY�ámo	"M5 �׃���ґ'��T|^�$]f��׹/�3�P ���┧%(�E�*c[���A΂��ϩVy�LBB��ƈ{7b����,��~)p���ܯ�i�O���[���U=f�c��P�%S�f������%<�#��@��7�pk��K3��Y
��`+�8�d���
X5?W��Hu+�pM��>T��	�X�F%�UBӂ-tu�����*�M)����Z����k8�(o4Q];���������j/��A��
�+��b���
���rj�}�ȧmK���wP�|�ph^��o[-9�B,�|�8�\���?�P�cѧZ��4@�,��7���i�05{��%Vk|���~�D���&cpM��~gBQ�%�F;�N�1�?J��⮆�U|�A��[�\�aOӿ�C�3�$E��@7N����~��u3�r "����C}.�����������6J*o�
v{
�K/��z����˵v��Ϟ�����C6������12*Y<^�,$�w5H6��L�b�	��6�D��h��%����U�����UQ])�N�I�����:=1�4M;�Ύꪪ>A*�!��Nߪ�$w=p�H���MI揷��a�q�q��Wķ4���nߛe扵覟&��.$l��:�W���W��0����@4�B�
@�2���.�7�+���O_��3Y̋�����b�]m1n���l����a���w���,�~;�9Z��g��H�ga2V��\ON��o���׆�����>
�F#��i�u�_�-ądؓE�PM��Ҽ@�$HJ���\8&�a��o�9�NrJ��zk��<	�r]���m�
���Ɨ mǫx[�*v϶�JU~b������>�сC%u[w��H��>.��EU��Ƌ�F4T�������,�=q5��gl`q��r�
��������k�	�y=.*D�^����wnI�) B��\ʑ �&@�.�+��*��	�Yp>�G6�捁�7��4;8��h:��cK$jj���Rh;�c�͐gΝ�M�}�#T �R�a��:ȳ��YC��v}-���~|�����?z��H���a'�;�ɷf���,NQ��^>���\h�f���i�3��:���T���E�-�J��L��(�]�6'0/���#W��)'P��)&�"]�EEMm�x�����v�ۮ���=�������,(�h%կ�(�ij���'a�=��g���@Y�LR��0��u���`�~���-��&I���;���m���
j���j��V���Ĩyej���r�u�L~�%��	�6�:�I�O_7�S�nc ���>�B�e���\�,�p;�4�(�"w҃ٗ�y?&EU�S=���J@^��B���l�� /pUM6F?�	o��6�A�d!s��JE������^ �.E�#E�����ВI�~���*H
@�rF��;��bb�?��>H���
�C�;9��bsk�	t�g�B�����x=�8\�%D*������d���e���-v��f�T������@RY�2�<V&@y�U��S��+�Eֿ*@�W��T� �]Y�(�w�u�1��0�&�&h�P������y��*tjs;����t���UpS ��BpA
)1�?Zb�Atn���F%��i%�G�J�̺�CY:���s� �n�s6��o��l�p��?q]��Z�=`��tN�u�I.�ǬA�"J��SaN����x�z�=Bᨣ��}�ج�����\1B!�jވ*l��CN��F�l,X���/�,=��;�H�yG�~�_`2ԛG��yv�N8U�Ty�Ca�$F�Q�B��J�uš�.���#�eu�Q��FD�m_h���3M�j��2N>�+��e��RZ�`�q"��G�$K����5�j�c�
9���~/ӏ<�	-]wZTP5����� �[m�$?� �y��d{y�E�k�N�Ҝ�0�wJ���ħ����bs��(���gv��{�!v�Zĳ�V��ǿB)ehJg�G�u� �e��	�˂9#,�϶Yz-��<PUX�b�1"�ޙ �h_��a^����}�=�0�X<�=���������p��et��|		S�x#��tH�yA�f�l�$}E�!7���*}O���FRy��اހ�4C��a�C/Lx�]�{�Z�-�؇��n���+�F�4�ɌM���NǃX�]��h��_�(Q��k��w{�0"Պ��R`�k����v�Ԝ'�;G�p��y|s2u�?ٸ$�����݀@��kt�S�H]���;��Wd�>���7��Y��g��.�?� /�lJ��x��:�]
5�+�yQl3���ܙ�	!���pT��b�v��V��(~9�D=25�Ȅ�U_44%w�*�5+O
�� 
��b+��8��N��8T�%�6�F�rn�]�o��)���7m3��ȟ��WN�M�(O�8��Kt{1Y-��،G�=n�r����A�����E���PEG�&Aw9�H/I&�ȓ�!����:�S߆B�^tM�7�Ql{-$#xhٛR���[+�GW�	C4�C�:-��DOJ�9�Ӽ�*t��ǂ��T�7��F�YRn�c������x��"'E|%�C[�a����u��ͅՙU\�Z�8��̚�h	�m4m\�^L��e��jo���('�*'b����ϊ�=�zHpk�xD��l�E�`$�xt�wIyZ��bn:X�������rP�7��ȑR;=��p��ɳ�G��Q6J�6�<�@��3/���Ĕ=��w"��PW�-|-f�u�� ��aaV���eg����@It#��͘�Gq�B�@��v���}��hv�>m�s�\<�M�����܌�q���%�J�ή(}��K��A�[�X���?e�k��:(��&�؝I-�7���sY���%�JJ�:,u�����'�_'
sٱ��`����X>�U�k �jn�EuE4���ګ�+�ϷϑG����dnRm�I��	��J� �M�.W� `���]-�_Ecv��%?(V�ό�����b_��X&��k��,�2��
�����G�󾚔K���ɲڹojtn�r-=�dxʍԷ)����9)�y6��y`Ojh��G��]o7siO{�~�7b��JD�X�1��)�����10�0݈�o�t�Ё�9,t���<��0�Sж9�����:�bs�<Q���*�(�<{������=�B��`E��.����T���n�F?z`��!/�a5�?��n��<��n�m,�Ie���7l��c�aqaI����:in*G�M�!r�Gyr��h���b�������$��A{3�w�4rzo��WBaE� O��4XM��z��j�����t��Y��lp	6��̅�V)�#e�t��;L;��=Hzoƭ��;*�;�U`�󤼩&�Lʣ~/�W��pY�M�j2�� }�7yZ���)R8I��Y�������kԞ~lc�̸��[}kY�1p`1A�-��AC�5�D0[�
@N�%�Z��F)Z&8+}�oH��`�Ǒ<k�D0H�?UȐ�:��%FV��!�`�B��ƢGn[7U��*g��|y�tx��K�4b�6ʆj����r���Ӻd���FH�M+0'_�PAN�x:�r�S1�|F��>�*"��Hwc���e�ֽ��\��+��tw��N��R�c���g���t(5��O5[ȵ�iS[��^n�r�y����"-�i����ݘ�t-$p5w}��k�v�������xibx�U23���AX�o�Ğ��Y^�K���LYe@V鸅m ���'�H�\"�߱�����$R9�R�z^�!l��s�K��p�j)|Lͳ�7��2_�e����
��G���]M��g3+����)]�Tpbu�!��^�OT��?ɗ��$������I�+=<��Jcz�(��y����4=��{:0�@�!z�6�,|u�󊭾��C��]e��^����c9�j"m�0x�Q��`O'�y/K�q�:�]e"���#��������ǀ��M�Sk�q+s�c{Q�bv�=��I�6T{ӹ~���[u��G�L�6>@�Y��"��M�;�f�3���W^���~}V���?��>+�ٓ5.7�Hy,@%y�2WAV��wXJ��g�Ip��5c'�B�:S�˭1P�.li�_9�!���R�p�u��;�������+��Ïׂ�����9
-B^F[y�J@w t;k��?���A���q�zS`�Y�)l��.moZ�cOQUӯ+�+�x1��s�a���ɞ�䂖`2�ф��`�m�=w���tB�ZP�6�F�ɻX����K���-c�����3 �S
Ϛp���p=�ŋ�*�U��1l�{tj5ݑ������:�I\p��<��Ys�=V�$������G��Ѳ��^��O��C���V?��r� :���đk�q�.c]�5���{���]13�\��0���i��=U?Wz��o�q2�'�36%]��f3%��IJ-yVp*{rvXM���岪�
�6h�}�)�]4�:�WLM �F��>����S�wGO������2>�7 ���L�S����x���Y�~���c��~�:�'� ��� ��F\��m�TT?��϶���$�Ƕ{�\�z�![�`��9���2�'&y�lO��#����A(;��-����$B]���# ���%�G��	T�!��n6�[	?�ӝ�5-ˉR+���X��.C���?�2�?΃$T
HI�o�,jYP��w�񃄒{����0�p2ImJ@�끏n�kd��ܰ"���<#�����-���\���?dn�P�܂��+D�̠�;�#�i����~'�}D�_[����=�j3� A�/��f9	������.Ç�9ϵ0�R�G戤��W��r�B=q�4�L��}TQ��[��Q����(e����H�t��U���W����p��W��Mя*%���?��X���K���cGIcи��曥C�=*a�[fp�!��|�O*�[eJ"�7�x,��L ~u���Z����(���N�|��53Ufi��x}o3<3�����ƌsD+�����#RS`Y�I�95�Q�M*��6+'�'@b\+Ur��P�O�T�p+N���-�i<��I���t�'�m�2��Lw�|���x�g)֘gZ�u���<ݲ3=u�o��䩮�YS	��un!�::��!A5�!z�ŠBz�i����,^lQw|�W�Q ')F�p�U�N��j�J.�Y����I�H�,�:�J+�<\Ǹ�>����и˾J:m��2�pr)4�>��0fW[d�t�96���z�3�\@���g�������_�Zmu�#���-�U!�a��� &Z׳��,�4^�-i��sh����Tj����~�)�]5�xp<\���>�`�xۢԖ���%;=��h��ݐ��x�8�$-D�9�Fj���m�j�"�#W#e���%kSU��Y[����+GP�V��%�uz����Z}.A���$H��㷖+�C5ü�A6��&5�,�ï,	���i�UϾ�֨��w�a|�c&T>�ť����'�8�u�}vtu��d<��+=O<�V"6i���}�/x)�*�>[�$�������^���J��v]b�p����L��J��38���w�iY������H�kgJ�{T�V�F[
z@Oo'6�h�MaɇVV	fr+���)Vm	h�2]����٣p�/�ur�vi����F��/ëصɤ��rz�M�A�G�����M+Λ���r�L�}Y����V�d�ž�r��~��}��s��QPu95�[�*��+��q�>��m���B	�!@�̌���4Z�y�����n�(�[�-YH��-I	��t����Z���_�I�*#/_w�8��S]���� &�=	��v3f�)_|2�/��z�,"�b'�{����"��s��VjA����p�YQY�q�\��٨ˆH�	
��G�I.��C�#����e�D�y�I.��}gN��ۃ.�݁�vr� VC����J������N@�(�1��S�/\Gӿ��jo]D�TH��`�q�p��ʟ�O_�dQ8�b��P� ��@��K9f��������,��C�ߘp<h���i����h8!6��iW8A�3�J�D9,��	�T��/�L�K�sG\��ﵝ�T1�Mv�T{P;��R�t�a���r�����S��{�K�lhk��d�W�h�F�BZ��l,(�a��T8�>%�چU%ܒ���K���"wEu�FDf�s�N+��}��!���gT@����?v�\S�����&p��"g�@�j\R����d2�˔�j�{�%j(�'%��ٯ>P�6�0��L-��0�+��^�8,��7��D���II�f;,ƟvxאY���Ӂ�A��˱z�zt���v������;��4
Q� �6(+^=p|�+z$�[2��m�vी��߽
5"�@��b��G�j����:�A�M�#O�.DB/�ӗ����BbTgyY�doaA�}Vء����F���?�ρ��	3�:l�1M[�ȹM!@�xP����2Ր���ț�yت;ٮ8#4Y����O>��(P�
K6���ίQ���FA&���t����o�x�Ó*�.n�"�e���5��}���)s 1�~^R�����;˚+ŁÐ�/(�d�έ���(���UNA$��\��||��<�eG�Wm�;���k9ͼ$�q�V�p:TF��F�����ƺ�J�ƅ����̂�=��-�,$5���O�4m��Q�L���k��^�u��rK-v�ؙ�����7���/B'��f��&:�-�Ʋ���RJ�*�F�v1�J��5����{��T	��X:�~�ᯛ{W�bM�����W�.cMG�6A�%�##�:]�.%@��߭�)�ɼ�7�� ��1ݥ|Zs{�ÇD�:Q��kn�����K7���M�����4��Jl}���!�~S����<H|��煱HT�^��7a��+���Uػ6^]�ʃ?ܲ�)�Z�#��Y~_�'Ia�b��a����I�5��f5,Qu��:��p�wV-y�0^@�bc�k��?0v{�F?Jv��؆���K3��u�P��}ȼ�.+�{�lK(K��W���v�%�M�ǞDwC#�7_��0��Ǘ	z����9�`��/�Y�s�u=����=N_���.�<ź��^�����2	? 膵�B oL��.�^���cu�d�d��d�M(��L��!�.�m*�-,��!b��(ϒ|����He?�� 3�_���_K^�o9=2��a�l?��e(��$㾷2U	�ӌR��ļ��׸N�vD �6k
��'�cw�E��+1U��je�qx�U/��H3�J��)�m�c���{��lY���z�ǽ#-���Ēk��w�
�9#�s����yآ*eO���(=t�Gƻ}�_h�Z;��ǽ�~UZ���k���%L=U��v�ز>�@"�nҶQ��|����N�T"���4�eݖnU~�Dӡ�u.4b� ���/�`����羢��PA��J���;xܻ�,�i|��9#i�{h����L�k=����?J�&S��à�G���N���	A=���s����{��+���8��ts.�u�v1�?�7��pBL�vM�q����m�}�N$je�u���t&��e�b{�s�5���Md��A�eҡ&mOsH��?S)G�u:F�78ݢ�����s݋0#"�����Y���Z�3U��� �)�և-~�,:m��f!�>��¬��{B��`UJ�A� \wp���m���P��%Ox(Y������]O�5i~m�������5�(L�mo8e}�>$b�G��d�x� ��BY�֗*���_Ʃ��Y\Z��;(M�Z�1+�6��B�Ώ0��K�/�v�,A��^_���"|ϣgc�X�r���_u��tô�����Cr�������qE�y�0nx�U��R��z-��pS�E#����.�7HU(��ɮ�p-ׅ���\���_F�,Ltu�6��	�F#p���l(�O�krJ���i���s �4��n<��T��Ʊ!\E�a d���a?ڔm���M�E��q�H�݂�x4��O�h���Q�Ք�0f�H�V0�ؿ�␉��Ÿ,�I�+|��a��R��!���R?�&V�q�h̟�வ�`�Hp�J�޷C�5�Y0�5�&��$4z�}j����J.U{ּ��$�o���'��p V��F�� X�M`s�y��	��&p���N�f��i[|�'Fs/Gj%=��`CP]?&��v���&%����%=�q��pL������R6DHA���3߸u�&���^�R\�<�"� $뫭n�10��X�����+��d�<���]�:?�F�|ܣ�Wl��<#4�W�_,@YӺ	)m�^�O���8�����$V<n�	��W��Y5,���Jm�Z4�M������JQ��(�g������šZ��
0�EXU���7���@?9NGլ=�$h��
��Q��*�GMJwD[�v�C��R���]s�7��K(x\��P��l3vf^m�+[��W��t�����2��ڿ�.���N���iY&��Ӽ���o���
����!N1��ޝ���F��eE��[:�c�
��Dz %�~t��5��-�k�YAͶ"+��|f�$��q�pX��D�G�A)��䕹��E�;o��Y��~j<���z\�y�����K r`���n�����H9~ƴiP���6��;�֥2����̕�K2-�r8(f��ck'�\Xj��Z��������oS�圜��"��L�j�^�h���A��;>�������C�k��-�����	ʘp'���[O����>�m�#E��{toJ �IW{ȷ�ۂ���v��1w\�O&_�12bM��f�b����+������,��|7Cx	�en���y4ڵ����m@q�"t������w�c*�¹�V5��3N��q˃h�Z�.=��!M��I�Qv���}|x+�?��VU�
^��:�r�a��՟�)���2D��f�P����݆A�2Ix���4����D𱵐|�r��<��,J^B�gw���i�:E�YVa#ާ���w&�L�!Q���F��x�d/ӼdW�Hs�� ��9mc�DLt�g�	mw]���`Z�OY;���s �������i��[AX����sx�z`�$���%B����D�YA����C��С;&$�y�6T?Q�'�g�������i��PoY�,$Hf�̕��Y$[,�KмŸΗ���lzb��K�$���8�kCsg���War	B�WQ�\죈$t�~��&Eճk롷\$��r��(�YN������~�>��5uu2p[���M�!�C1P];&5�2���z!;8��^�X@_A��ZQo`9؛Q4aC�j7����#������z��"����Dx�~�HC&�p�hut_����~k�74�7�잾��$p�g��\�U���ك.�Yé����A��Y-��W�-l���e���d'Lɡ������E 7��)};�B��2�)*��A�ǚQ6��&��������*�)���F�\�G��,.q�F�*:�t��a>�P��E&�(�;KX579Qc͚���u��i#��o��$��:�ـ�"o�g��� ��&�6�
�Ŵ��gJ���X?�	�l�����(VQ�E��Ds��eswCD�^�4��1��>t��3|�*�O*ԯ:)�+����� _��5*���mk�ҸvE敋sL�[T!�쐩��}soH\ꂠ4*1�>��2�K_.����T�a����ꙋ�K*�^O�� !D��\>�˝ x����F�1:NN�mI�>����}�YH��b�c�۴��ƃ9ȋBD���?HW�,�؀Z����_�`ߋ��(�_l�(0:�]v�{N۶�B*NF��ޢv��m"HN���;kF��I�e����|�&Usb�)��Δ�T茗�5'�e�G�:k�?6�
k� W��Xɭ
��ޮ/��en���N2���y��0��;~��RS�M��U�b��oV|�����W���\`���t�,M����x�<�n`�l�n(P�W�.-w��`�d1��U4���b�?�b�f#��&0��_Ԓ��Z3�<ܠ�W���ON��x�N8�#��OOW,1%�wE��i�i*\ػ�V�Ը/2�]q���Ed�������{J/;���n�h�H�
�6#i��.�9g^	ZE\��燲PJ�H�2�)3�'��k��E<*'�J����C1��s��*�I��d|4���k��?�BA.R��ԋ�0ZL.�W��K/����˖�ҮW��v۩Ď��甀7��V��I���ҀT��KN��AI�]�}ū�B�	�8��S�OL�+Ku.c^�5־99\���C������Lc����"ٜ�"���'6��G�=����ԗFk�諾����e��Z�Q^t��a���΀8?ɩ��˪���+E�[���R���(��v�9���!�@-п��pTSrB�l��%?�jv(��b�W�;��TT����	,;��� H��jI����ר� ���8=G:��H���(�*��5�B�+�.�.qT��J����/}Kp:\�Ԩ�!��;J�3��g	�菉n������d]l��=|��ż��ey������X�7��w&�9���^��6�u�I}���?�����aC����	��^���~l��
Ķi��-Qu�Q�u��tM����ַ:ZCe�u��S�+�<����T;��i��w���ðkwX5���U���K%�֠.18u����=D���f�4͇��j4���V l�R����L�Qߋm*�mu0�O+�ߚO��-���ذC��`9�Ӭ;_�Pz�4�y$�����b[\�y���9
� p�y�e��jE�k�p�*	MbDkS��"�������!1�I> �ANce���D���,y,h��O_(�[�+��\YUx>n��W�6����{fm�RxqΕ"`��$��v!j5�bR�^I\,x��^�c�4N�'��irrB���,+U�^�?n�X��E�T7�t����m߀��2�DXZ�c���ibu`y��_ñ4q� �x]1���yd�{�h3�_I� !�w8r�U���$��[ѭ������#�TL���Ai�V�Z{Z���	Y֯	6,5��*y�A����bV������8L+m-�:w��r:`JB���	�O
H���>���eر���z��c�V�P|:�ol�Gg�M�Y<�@�Z�I@�aT�&,��Go�Ƥ�P|�E� �$�F���[�"�|�z�j��`����Vf �uv�_��`ԏ���u�
����%'��,���,�V��[�N�#52J������u���ʀ�+6i�c�J��Vtu�!�8#x�J�}Ɇ�
�X�iL������H���d��cvZ�y`Y�=O	jJJ��IW�H;�!�Z��q�*����H[��&�fx}��v!ظ�ã�t8!G��N�dU	\����.Z0)j�c���.@��z�d	��ِ�rC�>&O"�]�D��敤6m�*��[+"��gQ<�N�s�1�BO����~�yϹ�Nʉ:��4qv�-Yq��N��Z��lYE��������^��F�/S$C�T|�f�~&/b ��u�I�CC�=g�I�敬
�tZ�T�62f�L�	�FSLKc\]"�F]�&�[�K��5�o��RL�$�|��������-Ҡ�Đ�DA�w�z�dn�;9����2Jù�|�z���������!C�l�prZ�_��u�pi��/�c��d�2p�6�oO�o�l��nb�0}�}k�M�t��J�w�i�{�>���Ϻ����)N�� ��ﻺxb���M��I$���0�������#A�0�my���y.n�bt+-�����E�;~�D0vZ��k��T��$��^���q+��H�,j�` ����e��	o��p�{5#c�M�X�������K�@j��`!�՗B
�����#f�]}�w�M�8$�s�q��P��(���e���x�kzl����{����h$!L8���M�&����auY�+4��.����>���zi����k�0��f��z����7��f��AȜ�s~��Č�U��[9�������ҼGd�R';�����'2�k�Ϧ'�'�Lge�������2%�SR��P	K�8�����T9�8����`W���l<�xE=�����v�"��	h��v�D��#�v��x�Ò<�� Oұ�+*ҔxɌ������ܻ��@Uc�}ZQ��u������������a�9���/�&J�=o?D��u-\h�_��5J��^i�E�)ŵd##���J?Dn�,g�s|qs.%�>�[?��.��"����_�~a�[3�q���w�r����BX�,�SQ�����_m�̋!�e3c��e�OKTT燉��;�� i��� 0�^q!�0��ۧå���䉕����õ�0s�C��j���Ls����U7�t&I����ٖ��R��,2��.�9P��+K�v6���EP��T�%MT�WJ�i��.1�v�~?C���ʂf�rSj�)Q��ʀ̉�����_0���K�lk���F�	tw�z5�X��0:.�/O)3w!Ľ��Zg+�\*�J�t���(�����q��++EE����z����ǥ�p�ei�w���.�LęԌ���C=��>�d]KC󮣟���H�
g����S�:�y���GE�8�=��皤��#,xz�g2�@G�������AkWumN#���xC�6[,���23�qz�	L��93�Rb�!
M��%�63qj���"��L�!����q�&\���C�̛��"�8�F���`v��L��A��o�S��V�"��?��Au���Re*�²�P��ӕe5@K��i��A)S�&<8W?���7���·$��n�2��1_�{�(����)�gfMx�<+�XU5�X�R;g�n�#}a��|M�` b�B��v���j���Д.`�R0;�>yoՕT��?L�\3*6�>zmn��-�'��ǧ��U�8��B�P�����)��f��������%��l���k��4P��r��3 ��L �a��IjT8U���t_�<��
-��M�5��r/(�,Oͭ$��ɨ�	����"7� SB��V��Ϧ����|���x��.*�b�;���G��z�3,c�@�1�P���ϑ��;x{HG��_rbUM�zc�)j���iu�����/���7�Z��c���qЛ �;�k�&���ʞ��r�<��~ZK!g.��F�,)J��ק��)*n�)x	-�YN:C4#.�4q?+������.<:|w�dP�gÝu�毫�Q����lW��_Rұc8��Zh�hS?��~��#�<(�u���C!�q.ۏ�	��i
69Q����Ƥ��r$I׾e����$ECnP2�_Y`�o��V�l�$-��\�8\�1�z7���_�i�r+hdi>!j��~1����`
�.��}RI�V�H8/�uV�l�6�A+�9�Q��n������>�?����K�a�I�LX�,�eKf��u(��z��l���Wrub�����A�|���"ƴ2t,�1�MW�\~b�u�a"�s\�7+ו��Y�M�eI�ε�o�6@X�
���*<�е6��)��idZa�#��d�0Ov��c�õ&O3#���ty�ưV�A�&�.�#�nZb�����J4<t�+�.�(b��`�~'c����8�p��"�!{�GfkҀ�����{��E�>'��kş$-A|=���ӑPW���W��T\~�}�P�!RSJ#�.<͎6���my�It{���aY�?�,Yb=~5�J&���^�J��l\��g���$��o�-WE�Ԅ.���&sz�d���g-�M먕�z(JQ�.X�f4��]�8b-2B0W~D��S�b�t�t>%�����<����9Z�<�:3��pӼ�S�4��+�
ޙ#�����;�d�8���[�{yb�EP���.V�j^���m3����n��Ѵ�.��/�æ�6�\�u�����'�#ַ
�(諩����3Z����4���yiRC�n3�^)YD���Y<���s?�Ђf���&'�1cC��i��gg^�heJs�|Q~m�M���P2Z,Ȱ���&��H�e@c��a�z���*�S���GB8����+�"�LYl�t�J��x�w��L�V=�W��5{��xO6#�b?۠$�b+vZ���?�r�>��e�s�&@�=�r�~�>"	p���=�]��ns4:8�F4��%������_Ԃ����V�w��H�]V�̜��l���`�_>&�.bxN��$oe�OM�"+��h�}	`��N��T�����~�'�n[K���
jYr4�D�T#*VM�6��dC<̖2Z�`�p]Kjs������V��1��}[TM�2���y�l�~0#�L3T�m�Q��W���O�/Y�7��j�YE>�$&�/N'�}�?�� 4�a��rK��e���De�]�'Oe��'*��P@�Tĳ����-dw_��
��:i�\v4N�[�E�e#V1���c��G�!��
�M�N�|��\���\v�j/�=�)��%�v#��$��7cr�hڎ�0"���=����B�v�݀&��t�N�����E�1@���D;������h����bh ��2����s�r
�ব� F@��Њ�����(7�*
��y7ً�{fuN�FE�S���0�r{���'�vI �[���z�*�U�D�e�_���Ы�9W��_"aS����K�������9̝�~��{s�u� 4��ne��9ۂU�i]b2y)�d�l�����ɑ��ki#?�A���I�&�+Cu!格�;7�\�n���� 8�XF&�T-�����}L%�ȧ�J=up�!>8L2F��/�r�l���뺠��ٌaؿ٤9_C��K��|d���=��0%q
k^9P|��63ў�7U�� ]����i�X��2x՟����%V2�=�t
Y���~����{鳲4Z�k����Q��BN�f~s�{��G;������4��SƼ*�9���sXU�às�e3�Xn_�����̀������B��s�/��h��d��I�wY�.U���z�^�ʮ��ԁ �Q��ÊJ~ٱ��9�9=SB���LR���D��y�'�f4�ݓf���3��Db�:~�E �g��䕇E�y
k=�)�["|L�ިn�@����z��D@M�#����^D�m�?bB�w0W�C��ff���أD?�F�A����3{O�);�1�]�l�>[,=�Ƌ��4�g���鞸��U����{\$���8��d"ń`���j�ĉ^�z��B�-���gd��r��O3�0�kjD�J�k��B�D�٢}j9��. �Rx�����J$�ʎ���r�f�T�Q\p�e��
�u�8�+��i}�`��c���S�O���������� �l��E��(DU��ʹw9�rVa������h�НYJ܌m�'�����bH�.��]���w9�u8��M��ls�����5��� ���+�q��x��)]uK��?��o<�y ��ھ����{���tF���
j�P��`�͚�$�D��/g��Q�H�,�!��li��Uȡ��ݤ�gL�JZ������p��yɣ�4¸\q5�V��AӬ82G���>P����=bT�u�D`t*�q,T����ۧ1e���\��{!����C �B&ވ�4$�װZ��6>��vȴ�Yt�l3�27��
�ņ�����(�V�8ά��e`�j���`�!�D<����~Z�l�XTT�y٢�VL���.��m��*fd�h������K�8g�it�e�NN��˥������EBl.���<|�e��nQ���I�݃�9���3��ߊTr�����������$DC#L�a�O�\J
��Z����dЪ�>s��a�d�ّ|�$9�H�k�ŝ�^�[3$�?W��#c�A�=ʵ��	U���|�Xp1g��p�GJj��Wt?|%n~H����E���i����x���1�|��֙19�M73>�x3��ۑ
�=��I�iN۟6�|��d�	`�Q)�U����Z�<��W���~�z�SS���fO3p�.��s{�\�$�U�z��������0�*N�����F܅j����`9�wQeEg7vR)M���{F��|�YfC،<�0�ܢ�<ߋ]�%�qb��g�$��I;�4�@l���&�hc����EjF>1��Jm]t���E�S�����c�t�Ah?fp�ޟ�i���Mmҟu�@���E��,b�Oe���3�#������\GX�+�4Ŀ"0]�CR�YPq1��n���vG�o��t��?c� ��ӊbWOn���É%.W�'���ȴgm�
�-�@����Ə�s�����yu�+�/ő���xn&c1{����yǯX�-�g����S\K;��r#:�*�H��D��z�+����{��dl��0���o}X�����j��X6�6b����c�b�!�ľj��W���kU�<��W�5X�$J�p���i+�=S�D���E�jN�I41N����7�d̓�yo���VA�%«��ネ^��ܙ�J�G9��$x>i��T��VdIh����ܻ���s.av'K�@��Ưh"<�뷿{��6��CTl��-�/�Z꯰�����	?'a\s�JP�9u�F�O���DЧY���x;���@ ��h���$�V���_�P���Z�f��T(�e������g%��y����QP�`H9Z� �_�#�Z"��d'���?�Y��(4v�����~���/sW���fJ
91��;�q)nO?��uݐ`�Ԧ�m�E=�|��v��;G>/b@�	0.؆�o���{L3���c�����G+��ep3b�,�$l��P��G��y{����ru��v���cM�$x��f��ୃ|�)�����@�9�;°)	�0��A��yl"��$m�Da���F4j:��k�$�;�݋H��A�#ݫ�KV�?�0�Y��A
ZdO&�����Y�Vtԭ�����D���ᾙ+��^�|�����XRɅ�T�b�RY���eX�E��؇ع�K[g�)O8Ŗ2RyQ!-S�RD�|��Ň��3P��m?���}u�rEɯ��v��ݍ7$!�Q�W]�%z��p�^D��n�n��°X�7R��{������m���{�5C�!�'i�՝��[�RY3�d�=�oԍE�l�:=���_؈�K�{1�HR^\{�����U�Z�~x���&*x���٭QϤiƮ&���8��29��L�69L�RС��ضv+f0 ohk=ڍ�־UK!�G)�� y�kh�q�\�jב��Dv�~V�ͫ
l��.Z㑷��%&&�.Z�ӎ�����1�+\޽Y�$0�H�!��$��pK�A����r���r=!/�^L�E���}0;f����a�P;���@gE��gG庫��_�mf���~� ��l�$2�*{����"3��E�w�o+��5���} 2�5���a)��C�l0v'��Mi!�J\�f$~��b�͛F��ѵ4)�z���Έ�|�`5�%۫��07!l�˓��E�Vy�y��7�����`���O
��'x���&5W�P+I�z�1��� OwR�����!��uӻ�;���m����������5�]x��S�WX!h����fU.��e�_B�J^�G�vB;m_U�NY�BV��<,����ZD�����J��p�HN���1���៤��J=������1dY�
�R:�������֦h����ߘ��Q� 5p?U@$��L��/�u}c�c���:�e]RM.����I�h�� !OE Z��4cS�#�5D#���6x�Mt���mҞ��b����Đ6�!�Wb(��v�`�� �1�&�A�D+�s�S��Y!�c�!�2Z�q��+��,H<V������V�1�W*Q�#Y}��Q��?�2��p�̬S��{���L����e���Qΐ�(N-I�Ԥ�S|-�s���R*F��!! �A�R���,�Q���.�Uz�'iFK}�Փ/��g]�|���v}透DQj.��ak�U^z)�$c�ob}�)d\�3�p�c&V$߳ e�	a��&M��
����4�_L���(�J�Iޙ/g�" sd��N�	�� �p�@���J�tH/ �jid��bp����	v�zm�-'�ÊT�Uڭf�#ؤ@��f֣��Ͼ\�$T�_�m�Q�n	��}zJ���-�1H���C�0w���e!�߱�\ĴRj�Þ��`&e�u�d�w��H+U�比U�o:�-_�VU�����:�ؙ��	>.�V
��]�s^�U�ʝ�T��Y��!���:�̀��FN﨎�o}Px�G�p�<9lӏc���_4���[�s��Z��8���x�[�!�jX%����8h�z��kX�A����H��萲0G�l�BkYvX{���C���� ������ׁ���qⴑ��l�A·ϿE����)��.P�f�/�+�B�.?Ocl$Q�������3���!�e�M��7�Di�H)|�~���(�2��M]�(Z��-K�Ɠa#�I3vxϞT��U�<OA�;J��=H�d6�-Kz�g�*շUD|�0���B����Iv_I�ij(�O��v$��Z�?�끆���
��&�Y[W���`�aqGe����V�&�~�\�( Q��M�%a�?��y����?��Bg^�O��op���2��^튡ǌr�D�ru��ԅ�iq�0�����g��.0���z�>)h���f��X��TPQqg��3�)S�7Y���s?������O��X�wb�_�<I����Tls���d�C�W����s�Oj���RMk�r��N���ɨq��rI�S���5�*��sX�;2=��:[~jO�ji�D��f�nu�9-�Z�]�Zt��G
�.2��t0�A��3����,s�&d|>+G)�3�xaUƧi��o���0Fy�����G1�2��G&�*(H&.$|E;���[B"N򭰂gZ� ��tFe��r�j�@�l桼�]�Y%KIZ�B�Zu�?�j��EN�|}����v��P;�z�]��l�ܖG�|��ya��x��vti��o����߭�Q�����o��c���o'�^�2{��J���O����J��I?PO�]���z���m�����ŀ�Wjc���< 8f���^�rg�Tk��������%��A|�fM!�����7���9�b���ֿhc���>Ă�&d�w�-���ЪR-�F.)w�,�(��%�F9`��+ճuA�1�OC��h#�y$ڙ���)G�����z�v�D��9�b:8p��_�"Q�	^��7�o86w��#��y�V���ˊ��f�ңê�K ��A1�"�y��S��,H>_���퐻�����ש��R�H��o��1��7;�W4P���X� �y�q�h�[��$[E+ �'Cd�+�N6����?�,u�n���X������r�f�I�� Y�����ݜ�B�=��{��Z�2'OeEj<ʓɱ���YY�0�����V�f��˃&<�jpW6���۵��I]i�e���Z��ʣF�G���<\�^�:��z\�c��H�,zu"���z�s:cy��2Dm&������{�Q8����@9yt���שӼ���R8T;W�e|׫���K�#t
p s�X�!��/������/Y�(�E�z(���j�<^8�)<�{��5_���[a /pnK8�d����c��50�ˠ��s�9b�yʅq�⟩7)��lO?qh�3��;~�8���N�>^L�ڙ�rh���W�I]�{oI����W�tr&�-G1O^ #��X{�����;5$�֐z��$/EX�ͨ�e�:�U������)#����4�r��%t�]��=�������ĻL҆'Ps����,#�^�_�.sɖ�}���K
�$��Mi�vu��S��D��Mܴ�A�4��B�����Ⱥ���"7�mv��,go,�B݁�̵L��	_��+~/�W�%G�BYJ�H]h��O]�#+�]��hj�R.���5H���N�o�G�P��ۀ����a`Zؒ��r�Ix��/(�os�k����3�x2���9C@�ݚ��*��
�]#1:Hv� �ؽW�	�W�`�__p����h4Yκz�@�Zв&����^uy^��@)�N��UK1)-������ �X.w�gsP����T���4��wu�g�.���ҋ�J�P��?�k{ClIKb[��&^�0I*�n��F������Y�S9ޢ$Uf�L�������XF2��h-Z�.N�Ք���}˽���@pI$��P�Q�˿��䬪/�;���0m�q&���B�B�H�i
2ٙr��D&f�`��4-y�F!���g|�y�d����ֳo�Y�������T��2K���y��F[������ �����i�����5��c#{�� �$�-�uǲS|�yH?RZv&�iQ@F���j�f(��M���,������!C�jF�z���8(����.���5�5���n���WGm8�u'uv�j>m*�c� !#`�Dd�Mz��1�Fx���@` �NɅj��T�p ���7�޶���`_B%T�����[)<Bf�^gi\&:A�T%5�qU���S�cl6�3;%�z���?(��/�a��Jw���������-Hs'@��&�-�����=ݬ-�[�~D��h�#�wL�N'=o�2|"��?iX8X�X���E���d��������)$�r���pYs I���$}��>ZAy�}�3�
-�Z�1�B�p4D��1-�ڴ��g�p�pV��b4��U� -D�QͰ9�ky���.��EGJ�1���ٰ�r�}�H�B�#��뤦e
X�����d�/O���^MuZnb��ƚ%GR2I����`H^OHA�܉,o�Ӯ��m�5���Z�u��>؎u!.�$���9Çb�$��4c��۴rXjq3��&E�3X�SzA�(q�I�fd�C'ܱBj�� ���#|�,�3�E�Y'B��!x�0*��b���^��5�qQLy:��CJ5�1eb�����B��tH��i@�J��ױa�i�D�?��Nd6��#���<�oy4X�� ��\w/`C�{�-2|qa_%��Q+�}��ab|��z�)�)�������؍���S�������� ޔ�+P�^�8o����
.��~` ���Le�Rk�D��SN4�,�ȑ�#��c��Fi=Z���_~Bw~��> ��x�xgu@)zIy��TGT��Ov�Y�G��>W��#�����0��t�5r�>B�~C�dR����dO銋|�5��kzv�e��<�R5��r����?T�y�z��K�f��IY�e�+�;���	�6f_�-s�/���wL��!�oۣ�b�*�Lid#�P��F�n����l�W�{�rm=�D֕��L�ʍ��j:����S�芛�f�퍒��E�b�#�|�,�6m���z�%���ފg�y��V�����ӽ��;���.C�0j҆)��ar�X5����U����o�J��t��T�I���fa E�[ncr�̒ۛ��%�Ќr
m�I��UI�\F'������Uq�����b[>�%�x�����9qz	�c+���]}���g�SG���������1%��7K������<0������x��hŃE�٭@���L��rb+�KN���� �g1t�4ezl�b*H��O�mG`M�c�c�cup#2�S�2ߐ���А6�fY!V3��플'�b��Z����+�u�T&�wz�M���䜐G�eR��]	�zn��ܬ�_���ϻ4yt�1:�~
N�8�μ��	Ly��$([�h B��wtxm�1,2�Hc�P�	�=�.�7���&ۥ駧��K� �@�GN	�;�lk�)|ХB
ѩ�j��v�}�S |E�ȧ�K���Wf�|��'���D.쀙����rXJ��<�o�]��Cַ�r�E	����&��@G[b;��v�A�3l��Y�m�N�q�9� ba��c�WM	�H��k~r#����3RY'I����X�!S���'$Ƥ���WM���.F�q|�z�q\�4��K;P��MC�:
t�.���2�x&�'%��@Y�ỳN�J�e���ql&�ƞAk)�L��K�S
��	�g�K~_��h#�A$6#��7r|2�]\wNىAp����NxI_��,I�!��
h�������czj�����_�0Z�K���_C�2���S�΀ds�Eh7O�hd�C�)�]�3~;:��z�)��S�����75�|�)�,��h�˞�\wu�{�/���:�D崔�<���R�+P��>?.�;���h�Ȁ�:-r�1^�ă��(AJ�5½�*Z(4�t(�Dj��a��O&R[�6w�"1���ᬎ#5���_�JcB_��Rog!�������^f���$'�����c��9t�@X����1�=�Uycf�
��~,�ew��Yj�s���	iyކ� ��E0#Q9a�ӋdOT�D���Sa��us�X����(>���������I�?W�	͒�tD��t�M7u3 m���v�E��j~�{K�G�u�S�gQ����X�x���	�M����5[��B�+�ш���;Mz�k�,?�T���)-=�])���OؐʽgB�A���v�H�?^Z)A�͢����$u��Ur�NT^�C�bc�D�U$�v���d��@2Z���K�GQ��.�c���I%w5}Zɝ?�7�M�"B&b����g����U�O�SB�C -�*��$�C��L���Vs��ɫH$Ô7){{x�Ԉ;`�A��b\Zܗ���N����0����p
08��ȠR�h�`��������lȱo�9��~m"�JE���\ϫ>9����P~0���ˎ4좫�J�	��g���+Ρ��!KjA�<F��T���˲{��s�{��|������U��%W�C��j1��sʩ`��p��,�~b>_ѭ��c�mp	��o�Ѿ�Eup(KU�s�G]�Hۑv;�Ab����e1C2���t����s0NN0�������0?O�i�us=,Yc�xJ���4��� S�F�:  ��=�c��+�_��I���:�7�.5�&���ҟ�[&�\u�&�߿�$�\41�g��c�ڛ�y�1-���2���U�l#���YMh%�G�v�m|?�BM1h���oi�ǐ�H�z'�~a�d���N$F��
n�Ry����5����l(�)�:�=��O��Bo�\wf�j�9�Q����pE�u������kDq�S�U7����9?��^�xY͹%OaD�.b�Zd���I�_[�Qj*�l��r#}�F뷈�J�J�c�7_���d����[o0��ܛb�c}p��>�ڥ�o(}�Kj(bfKRȢ���CT�L��]Fw �#���s2]o��҈O��Sk�� #�"m�2��!�����h�,��[P�N\����]�gO���u{��3�x�����A.sKM�r�!Ӧ2`ϝ���k3�9 �~���yP�o@�-�rc���9!���}���'6��X�sn�{3<���+$Tq��SD` ����~^�����9��r$	5�دJՊ��cA�����8��8]0�8N����;Zf��PMl(T��H�G�����S�(�q�R��T�9�w��0ߖ�4>��G��D�/g4T�|����%� 6������5Ʃ	Qf��hR͟I���G��W��w�J?A��gzΩ_.u�@?�mn�U���~��?�MF,��2,~(x�5kj��˫�p�x�LG�� �f��u׃v��}���ɔ��~��o��>�c+�&�n��WRh~�琁���^�eV�S%����?� ���u�D~�^r�7<�I��o�MF؄r����@pA�ϵ�7d�r9���5ݕ%���8yȗ���� �4�,>��ᴆ͘�g�5n�m�����5KX
�����՜u�fa����/�,�� �%dx�m������P���{�+y�HE�D�+mř�s���U����]mv@���oMZ�|T?9��/7��pv3K�tEN��T�'Y���`w�@)���r��SMF	Lu��w�0ێ �y��^
o�.�v��pr)}�|��<�{�� ����"��Iʮ#�[�@;π�3�)�bڍ���G����R�^#�Bo�@����_��(w����.�kW����*��nd�2��_����=ڡ�j���d��=;�G hI��/U;��&�[�}�~y��5=4��Z�h������R:�A��2�s��>8{�Vo1kM�G�W�&����v(���i���/\�4L[]?�X70�e:�,o�睧'�Tg����>�S:��l�nX��R����(�&��j%7�~t�W�s(2��(���7S��w�ل>͈Lö��y S��l��֍.���H����gF�&ĵ����U�Z�c�g"}�~��(e:����p^��&�8!w�i�<�!���pُ'���=�CsТ/�nn
�{� p�Ē�Vs���6k��	�~�V�ѽAea����,͠6DT�'��#�Ry<V���JA 2����m����AWg|������+iO���pg��0�a�Ș����c`̼�yO<i���o�����H��]��g��y/r�O�)�`F��7�%'Z��mT�^�3-��T���`|@o�����~�O��w�8=��;�g�0�>u_S��W�4"l#,ŠF�4�`��/�&�	@dm���L�^�ci!ϺX���
������`�P%%�֤��]t,j#N�Y��)��a�.K���C$d����{Y�eOse�����`�x���!8;��x�Q�m�@�G�*�����`�s����h1���AI���v\3hD����R���*�|��ƫ�Y1@��u%��6V.��{=Wn�H��J(��jw�����Yyq>9�
��d���&8��RI�9��V��Ϸ`�$(&�Ad��Z�pk�nՇ�K��[W����~d$��H���<�<v]�]�+W�rC{�J�_�g�0�N���HS[(36W�5�1�B��`i��~	�����Η�y�	��#��6��pa
�ʫ������u���4��4	-��_D�(%�\�.cV�蕠��	�<�4�9�{e�	�X�S���ׅ�󷍶��O���;�@P�W��W�N����[��s̬��@o�s^�����N\H4��f��ER1~h�9C���Ir��ۇ�({S�#��Gbu/el��������,�sD5�����z�1��`�FL3u�ZV%$����[�*�uMh�%X:!A���u�k4l�F���בr��� T�>Ufڶ��w�q,�ҧ�NS���{y��V�\1]"��Ɵ�E��};΄�P�G�Y�˜j̩�OD����v�`!�,�n�<!�����������C�:|��O�9��;62�f�@�������H�x�0(��Ń���xߪ�K��Tm�����,W���}��n!�:��\x�����fwF s�f���5y������5���B�(��E�f��1�I�_W�ܦ�-ޚb����	�M���!#�E.}C��������8?*w�q󊽒VKZ�BՐ߮˗�C�����sSQ/X�e�Q�=���Y�Ə�B�`�RW/U��2���B��B0W!�4u/ k37��I�J�y'69;,q�!s�ED.6�e�U׻�dc7�o�6a�s&ZY��m�7���'�O#�Yb���;tZ*$��$�M�G���/�I1�8qu�]Z�)��k���P]�X��� �3��y]<��Pi�`� ��hn~�x�v�~,�����G�M,\*v)������~������V��+��=�����ս��Z�u�l�v+�T����:>�'tC�p����
�qwI�+6wӒI�s�k���?��x��Q����DZ���XG
�xp��Ї��Լ� �X�m-�2иBN���, e�,�sw��W�]�~�G�y�k�:0�k>B�H��؂4�����9��AbIk.e�����H/�̭�V��'�j��%��5f:Y9F/�;�aKU���v�7=Y�KE�.��9!��������h3{h	�uS�C��� gB�
�9�2�J1�;��{ä��Ժ�-Lݳ�˚j� �%n�����/� IC��y�\�*l/�X������{4n�v��q̈́F�y`� I���:����rL�Kq���(�!U�y&���@�����U�A�Ht�DykwK�Bx��#��=�+���!Sp@K�v$_
_�i��В�$��p]�m`.S�YƊݦIV�!l붿D~��N0у�hHTpBo�8�wpX Ž���#Q�MX}LI�$@�K~./�����C��ɞ�N|1���.�5��^��y�q�a��Z؅!���۰-I�Gs��܍�ď�cT�"ݭ:r=�x��m��n����KC3'�VJ����p�4Q(?Q4�Uc��l�!^��Ss�tF��7蜥���B��]F���1���T�T�	�ʲ�;D���D��p������O���<I����ͫWB�h>�,�}<�p�S48�?��}����~�*�˱d�Tĉi���^��۠�)_�Y�_���55cEa�	!i)�4���bq7BNuէ�T��ۂ� WCm����g�^Y��荶90D����I�_�i�"k�:o��sL�5`=6�JSGla��Ꙥ��N�h�Y�[�X�-�]�?��I�� 5��4�i��R@�����&�k�zl��>�ΡA�;=y@���,�x>�!i�9+�n|��Z<�@(�\�r��(��P�Eyi��	�~�ѭԧ�j��FB���@��*�RPi�J��dh���F,�sP���A!���e���i�a!���:��J�,.� �嵦*Y%�wl�WI~B���(�D���P69��cXj�79� 6�v'#B y}-i�Z���tr�p<�?�|֠;Я�Ѕ��C�+��9j���%q��f�cuX�&��[Ѱ�YG�T(���V����޵���0,5}c��5�c�v��œ/C�F��;�36e�ԌKiØ���+�����7���ب��\eAJ�5'\hE]]�Q������'�l��u��x�/\	�J�И�A�"��Ú/��>� a?g���y�W�/�hT�
��	mQ��z�CJ��T��	�h�8�C%�ػ��zׂ޳����SW�����.�����0�(���5�y�g�D�|u�"�~]N����gR���q���j��]e����,�Q~: 5�
��f��i um������|��1ᢦxi.Bn�q�E�*��^	�!+c��Br�Z̏�I�+��;Tq�5�o�jUjt8Pt��<����=��]7p~���u��J K��k�DC�[v��p�9X��&�2CLo�<�k�&NY�O0都 ��u��&Ʀ�!!<��/R�3i�+����)������@���ݱ�A��=np�-���ߋ�dI�m�<l{�/�9���8�&-�}2EC��j�2������K}�ۨ3+��t�_��>��4�*)�.vg��*v�->,½J$[�H����#|�~p._~ϡIJĖ�f��FbR!��y�{UD.nA�nJA�P,/��m�:V�}}�1a�=N;����x�'p.U
S��>\�Q���(��W��I�{�_�o���s��*�57{�f�yo�I��<��0AO\㗪����h#\�8��m����i�"���.���l�h��,枋 �x֙\nFxw�jr���,�D�Z�$Y���/=K���t"i�e��`�~B�զ33@��õ�����#�a;�ʆ��xJp5k�a���Jb�L�Z��j�;��q���=d��e@-����oc�G�j�)�!��[�_Q������_a��H܂�6L�hi���"�?�a������������cg2�lz�3[�}�i@;��E�g��$�'�~}I�u����	
S����^�V��ؤ�Wӭ�*[qK�(z��Q���(<���҄�����ߴ^W���&�4A�g5�fQeTMP�Uɲ���_�ׂ�#>e.!�J�!v^�<�bFݱ�B;�y�bί�c�)�~��l:�n���<ԔB.��Lyt��n�8�4��g��x<7y��Wx&��)��	�@qd���xY:vז�`w���~����>�)p��K	�D�/�H2!��u�'E�3�5�">�/��3�.��\hT�?b�w�f0~NI@VP����_�.w��Q��Cτ+Ux:m#<t\D�
�ت/������4���BШl݅�P���O��nMd���t��;�-%���}j�\=�
��%>�k9�|=��p0�7�~�'�R�n����=ڀjG�R^�
_1d�a���̮�*��������ob�
 0ܐ�L�;`Sd4	w��UXu_G��Ďyf��{�h�<"�}����a���\�[f܃#�iDH�kT�2� ~���
�4e��;T�l��kv4�lc����O2�I�����}�#�I�Iul)�IU~*���Z/�;!d��Z��n�8�ԡ��ỽ�� ��4�,��a�0�d��ߤ�~d�_p�᪲�-�ZT�е�u	�/a�yQ��r�	��ӛv(V��#�CN#*���Z�qd��uH~���.x+B��Œ�F��d�$ɿ�XRY��<�Xbͮ-�N\�n�k�6{ăP<P��V�$ٞo0�*�0u�>���c������B�xż��o���z���dr�D�SΙM}�~`Wa9��ĵByD����S�mI,��i�&]P>US���7-����� q�_.B�z�Ub0�������r�9L�{&�u�>PR<R$�jao�JcGW�KL��'��n#>��ι�>�����/��K��HX`���A��f9���n�1�7��D%�Ɣ;���Fk2��L��d�߽' b�[g�1%>J���UÏ�wɍ��2��_ 0��D��cc�?���j(��p�8�je^9ʈ���
�{�Qz5[G�W�>�����f�9���E���^�S�0ݶs���(�~�Œʣ��R�΍|�:�A�y��/)8��ǣ<��e�p�5U�6?'�)cB�/����&LIo�Y�Y�"C�÷��H��O��U��^��Q$cD�� ���6"��^���L��M�Wܧ̸;�����8%�Aϱ�~ۇ�U�^>D.&2 `E�4�[u�}[�%�s9��i(� �둏�_L����������_��c|%ˣ{�+-�RQi�}*ne������q�9o<��힞p����n�q,'u���%](>W7w��O�9��*�!@���Q����L��OK��yÔ.��F���Ok�ah|֕L�!����V0��Y�{(��o�A�#�L�s�6}�/�m&�AY�>�{��ل�����b1����ċ�2��}tJla�w�{�$�a��
�pТ�=���T�����;�%>s0�t˿�-�_#�im��jO��X��j0D2FAZ~@#�/�ׂ\��z�@��kX�yD�3.r��0x�^""�΄\���(�j4��*�,i ���سK��PD��C���oy���v�-�8��׶����|�[fm>:��
����.!����?%.B#�{����y�8��AN�A5�xW߰�/81�&vx�>��P`�����^�D���<�+b��?�3�g��m�^�L�,�S#?�P����x�;�kf�J�G������$w> ��:V�|
�M����!2�"�\��)����F�ִ��x�0"���ş	�m�D�|EQ���H9dU�FJ��W�:n�53[T㨸�<�];ycJ&稶�GQ�e����ҷ�q��u�o�5Y]���F5�BU�,�]6���n ���rd.ԘQ��]�֐/�qGT-rc��ZR<6m�
k���Y燥hD����F=y�0�IqLA�u\���h$�-��7���e�'�n����q�E�s(DpG1fn���7��w�)A�1Sݾ:���f	�;�c���*��u�x/z��Y��^F��@@�+\8���b���ߦl��Ԝ��=m�p�`���I�,�Sgp_>v)l�d~t�23k�p���T��y�["j	q%�'�ϱw|z���D�.q?b��Sx}N���r	�[T\����
������ ����"��#qV+�'��mpZ*���-�*���,e�J�pȔ&p�p�BRd��#����$~T(h�/`,����
�4z6Sv˂N�lכd\��o�8/�p2�[�bs������̞�,��S��Kj����õ̺S7��R-���X �S?ea��X�N�h���� ��H�s�8(;1���פ�UyZ`�XD�m��c���F��V�:�H���4*=��6��2��E�[5%�(��H���{����+(Vfɒ�t ^�����������4�\���-ӯ|V���1ڂq�fNm�X��p���6ҫV�Q�m4�`�C1T�б��ͫA:��|M����dƗ�+ ���E�`�+�o�ev%u ;���=�a�je&Jy�w2N�~�Y���@n�����<���K�c�IRI�S\�M�;a�Q>��������|�O��4u�Y���!W<D�v��{���~��I��;|�B-�qՂ���p�||c��c�;5�����>ɲ��xX�r�]�m�>=���w���Ji��4�:���Qi�fC��K��yh��*U�v��^�@Py�E�6�/��Z{��5����3��»�T X~�M�"���n���u
;��ؙ���)"k� �ślC3Z���7�GV���9�z~����d���G�����}�3&�|�q��To�Y�\��e���v�$K�c�r1��@�,y�woϬx�V��YM�K�١�4C=F���/(�نĿû��l���XP��4��䝹�կ�X��UkA0�?���K��e�u%��Z�-������ n�O~6yL{����h�&�quٍ��y�m�=�m��)�"������mjlV��6��ؓ�@�~�T�w�1���G�>�d��U��糇�o� $Π��6i��D��{�/6��M�oޟr�7��r`�d���V��4�4,�⌳�
>�e�^��cM�P�T.�7��4��'iy��!��5@���]/ˤ��l���v���8�� ��mT�dN(@��D?��^YP�VѶ��e<��z��}t���k�TRI��0�듷�cD+ϵ!���������,�vz�x���B�7���WJ� lA�ಹ�}t��&���'>�
�����������&ª
�U� sab�w⒂��O��Ȃ`�)�i{,��)-�o��a���q�L������w/Eh���1ݩӦ��d��_��|���_��ؔ�Ma\�B+�����q�"��O��V�����kX��Ա�8 �}���,�s03QI���`�۬���T5��J���+@
9^�rdk�Y�ztSPs9F	np<5�v�w1$kH܈x�e��Y��+��Y��f�T0��1��� �� l�;|�a����r�0	��z����D�s�ڔ13��l9��9�'���p�o���B�[�78��/�Wv������z��/6h��:�,�㍔HHc�EG��//�,#S/�6��8��y���`f���-�~�`O"cBBGȷD�����.����d\ 2�69u���d� �n���0X��u�z�VHې�PQ;�Y3�UQ�H$�]�*�M�H��2g.�p�IANM�����=|�pJ�'�a��Rc�$�xI�������r|��jO��q�@�@?۴��f�����.���S���nd�uZ��{����Ig��9�r�����@�����UUn�E�n^V�5Ş��/�x�&���������4ML�Iѩ�0�d��ul�W]�C�T,�ϒ\#,��p��啉�F͞���`j ��w�����/n]f:��}�>��m�	�G�ld��u>�^�=3���D���,J�4?��) c�I��V_��҈#�.h���V�B����l��X�	�#��adȦ$®"�f��uB��b������"�b���p��0�b�ޠh�7��2�6�S�z���N)�ӫ��#�&��U8aDe���<����]nzp��팾1������l�x��ᬰ=��*�}�����L�C�*wT�����//��A���A�f3$�]����865N̑�샢M�'�s.�T�-�M��{!�Y���&�.�����i$����d�Ck��*�w�;�,�8��"�B`1���@�Z5�
�]eۓ%>.G���a�Bk���N�-U��[��d^�ŝ樀��j�'.k�׶Rb�]\g~)Q�9A�^-Y�xK��U�� Ғ�g��kQ�4 ���xj5X *�K�U�0~� �;�
Rkxkf�G$�N�Uc����/�Z�QJУE�����m����cP�:�~E<v�|Q[l��5�5|&�kPM�[��OV�4m���q��i&
o�H�9����߫�]^�|Q}��&H�	0���u$9��i�(1�-�߈y���yMt:��~���}l,ҺU���%�q���'�l� Z���a��e����f8��U}��f�&>�0�Q�loX��W�BtT�{^�c������d�Q~C�>F�(/;Щ<y�Qm3���W
�S薨qk{%|��_���U&3$@$����7�GG��������#�jJ�V���P3�=J���[j��I�Xr�9�]�q��̀C�hE�%JR=�3�J���[��\U(Q� ���HzFX�¨b�̢]�$�Cۿ��~�UV�g�NmY~GRr�V�/4�k)i��V�$��J���X7��_�ů��Xn�E��ɵ���q�-09I�W~�T��AlHB��@�V�'���~��%�BC�H5@i��=�8r?�:%���*G����kcЎs�]]��y^d����P�4BcB��G�$�,��t�6L�N?I�e�|�6�@x{��K�A��"F>?�?��P�������C�&�.	��d��)Y�Yk�FX���y�ͪ�*���X���]��D�8# ��n��Iɔg�~[SJ����)[/T�Py�,��jz����}���R��#�vRˡ�J�&+K7 �a���l+D��`P�a�R����He��o�]8��%�p����������P>	�3o:'����}Y5�@b(ބ�i�xk�j�9 k9���d�K�&s���iL��$�o�]C�	���_�p�U)�!��O�r�H���qC8�M��3a��'��g*)(����r:V{��Z���o�r��4�83t��W��QPUnT�3�(�#C� ]���>�>�_&�H�{�}�ـ�e��a��Ñ�X�Gp�Z��C���A�a���L��@�*���ҧ̰ʔ�ݚ31(���u�L'e�]��=j_���Ar`���{�&�%�	c���I>����lmrN���e)��4�+�A5*�֡�"�~ GA$�`8�������u��z�yNc�*cA���Ώ��j,6���Y[m�)C�r���75����?�^&\��_lE����AB���ֆϼ+(S������6c5�a�Pޮ4����=?W[����>Ca?�5a��$ڠ> 9�շ.s%M���o�L�=.�~�T�O�T51F��[�Eo��A`����l^���Ʋ�ne\�/^�4,22���������ߙP��r�?�|�ei���u6�y�)xC�	�3��Y�d��k�]���_����^��S�#�ޛ��l3��6"��!��.&F��.�i���8ϗ�{�+n��ܤ�"V;5�0ͧ:
��� �yb�'���H�񏷲w:W�?�5��e[�h�������Q�Y6|%���N>x�v^=��f�\�&�jʉ��9Ɯ���Z�4AN^mn�]��vL�+܅�s/>Z���׺��mM\*EM����]Xz&g?��>�Cz���J��Q6*㙐b�D���l���fϯ�N^9���ӫ�un����-Z�fi@:�B�����_N���
��ڮ|�o��ۉ��G��2�F���7a�I8c��!�� �%T7v6y�Y�Q��h��{=�����'>�|�}w�x��x�rE�5&0������u5$��59��&�����S� ra��(U@����u.-����O1Q(�'/�*�
�hƜ;B�,0�E*������SU}e�:FҖ�)�AlY��}���{nq�s� J����˯���6Ћ�Ť5C�AU'�Č<�*[#��!2��ն���Q���^ָ"#��@R��V��c��Btx�	��ı����j��l��g���3�:_�H���������E�����ޱak?��_M�Ui�ߑ����#ƕ�G{�)�̍�D� Հ���%7؂�b��0	�b�H[���<%����T���.��`�N�B%Dqg�ڱ7�G���|����_�q�Q�l'��L^V�k@&��f�{�F�Ð�<�Ʉ��~�[S)>	&�4�M�l�:��6 � A�-Y��O��vD�^դn*�љF����P�z�8)đK��ѬLC�bK���_TY������cO��%�_����Bd>e��b¾�
5���gv�,[i��:<$7��0�`��^b�QUn7 \
KN�]�:3�&~�Wz6�Z�'}�w�}JHN�Y�����>W���5E�ЧV|�R'���;�s���Jw��Cꙥ%�M"��}"l�XG�K.*[k��O?�P�R;��&�.��3N��WI���r�gX�N����ŀ�@w�� Lӄ44��N��g��%1v���5`|F�z;��Q�8��ϒ��<
,����^��UP��~R���l�������w�y��F@��.�t�����YDiI6^��/f�ֆ�Fq|�|qq��KpҜ�jx�̨&�w>r�G������qD��⿗G���cJ���zo��`����H�4�E��~fzD�(I�?�z�Z��#��=��Lo�/(�f��n��ꏒ�cjn��hĂj<4�Kp�o7��'�����dW��L��w�9-�T(g��.C2�,�� �4�b	���Y)�_���6�%y���@C`�vI�������$[Yj������6L&��b��n\� ʫF�|*w��ʛ@����&��['W"�/��G�Z��E�U4��Ͻ�^��cJ� �Z�(�Ư����1ü��3��o U��W�{�S��L[������a�k_Bn�E�^���&����E�aw!Gt�`G��~B�ǻr��#]q^ME�;	�1���XJs��ƘD��B�eؐФ�r��o���>����o	���ur0;�M���������v� ������nM�CKSA��Ƴ��8
ٖ��v�x5����}�Wپ�';���vy+R��V��SFht�	� ���ih���8�L�Ӷ6�E���_��S�|�4}���A�*���"7�8��tƄ|���Бjt;]��R^���1R��N�^mVu�T`p;���ʑm_�B&��X�7�� d/s�,W$L���`z�շ�?i�!X�/�Ta}����hpIűK�^yFc���,���B0�35{"�fљ���IbLG��d������&�l�i��d��� sacE���:�&K���F�f8��m����]�=�\��'�N$`�"	�-�EӦ�^���� �8�Ї<��0���Qs#���"h��~����s"0���|�gw���r�����U�b��4)��	\����f���,���@�m^.�e���;<g9l{���o�'��DԺ��|�3(�2��A���dv���8�^@7dM���ӱ2#9�0H�=%Fs3��@�6G渕R����������x��իw�����1|#���n�r*|j%��o�h&����n��y$�MW����Í�C'�=�϶�����puc���Nffr�	����y�1:�̾]=3j�}6�AwQo�'X@�bݎ<֮�8��>��)#G3�Pu>�<I1I���n�e2�����ĳ5�)��ܕ�}�SF�m	ȵ�|�e�v�`Ot��/�����6��p�{W����������|@Yy�_Y�)�X�U���&k��sh����Z� �k���
���'�"�l�P���7eS��3��[ߘ���� mJ2��-��t���y��3��������ק�.v��-�ᜊ�*�:��c�T���1���=�Y�TkN�[�)�n�)6���o]\YH��S���4��"��
�N���xrْ��G$��.��6`R:�U��K�1�-#��Z��C��|5B��d���Y�s�7�d_�ŃpL~gD��R�ٲ�����=���U��M�f=�Ҧ����n�j��AB�G���� Q� ~f�X�Ap�y��<�^���s��pJ�_�<�£F�Z��"���W@(��]gK��#�<��H' =��>b��2-�?�ۣ���s"��ħ�)�:��SǛ!��qA����ܔPu�$�J~|�W�r_!G��J��R��R"7$u���gWY�{{2&�c�?q?�jr<�a�&"����]�U��l�x�l�m'B���ԗ���i�����5�����M�6��y�&9��U"�l�yd9v�l�����F]g��Ґ�t�L��X���=���"��M�^ܑ�=�r�;��{�ҕ����K��?��P�O�ͻ��-
X��dA�v�����u���H6��ّg��LD۷j`�&A�E�.��@��|�%Qiu��!�:��o�#`dH��}k�L�9"���ǽ�1��N��M��GkB��B�]�4��'��ݳa �r*�6��iC���� SFe.���͙Z[�Oy2:^m�z��%X��6:z���;��k���C���z�����>3�xMi�' ��z;{��d(K�������4�~e���,>�S,�Q�u�oĲZ�L1��mŜ�FX{���f�rU�LQ1��]���xN�PO�WZ���s�Yg4wrj�2s����]<I9������Vpfl�v�C��
����W���D �����:��=��s��qo~6l�\% �Ӷ�>��T3i&��	g�F�1�G�T����� .����mC�S��1�}�b�?0����2���b�H�G�+�H���=��s�h���^^>��,̨)F��s=8k t�rx��Xqa`��{|N�*fj���h���]uq�Ob�UpR���mBF�.�v!��SS1�3��ֶ6��1A�A� ���?�C�h�	�J�E����R	�ZJ��S�V�mJˤ������^�Y8t�܋#�k�y [W��,��<�4���˙;��S� �­�?�H�H<�e�Z��KA&��|���TJ���aR�]yc�!�O%K��-��'۳)�(
_��b@�]6df��,#�b�����@0�W�cܴ5>�6�J����@V�+�v�E�ys'"R�O�	v������6�p }���֧���ﾠ@,%ZX;�,�O9-�22��=���gH^^������*���t_C�r�0�5�`������}��eT��ku�qݼ������0�㣰�B��3\V��}�qwI�R��.~X�r��u�4.:�C��V�sq�;�+�zp`$��=�Z�_�N �>
v�~Utqd�\:J��u��C���6w��&�/eQӁ�ҧ<Mm&_@4x��iC�u��y�m%D$���&��G��۝���3<l=ֿ[A�~�Mt��%B6E s
Ƞ~BK!��#"�wu���bز9�/�i��T$Ӵ���N���8!aOߨR.Tl�DCc�B��Ѣ��Lzӫ���ΣA�B:��>�u�Q<�T[-r�E3 t��n�S��<c>�W��n�O$4�*�a�X��	�D�u�:FGSM��2@,u��,��}3��k#�ݗ(g��_T~�-��\��F�����i'��#�����J@1e��J�i�%ض��%/�82A���8��,�1�[������z8	���V���BT
=��$U�<R4�y��� �	�~�b���gM���T���wz�A]���i��ҍ� ��Ss�/�< uå$lT�:Y��A^ljsw���1����}�ԏZ��d��|�	g��<�p- ��m���H��{��ҍq�t&���t��"�Ν��TEh�ֶa��3G@ea������d�!��/�		��x������0�
~J�z�y�%}Aj��"�Bx��E-�D/�'DY�{,BG4w�/|���_pN��g�zx�Xyf3gE�����R��^H��U��:���3�A�=�a/_�H�d��f�J�)�ο�� �$R�^Z��l�R^��!Gn�����\+eQ\�y()�U���Zw����L �{i�0��L��C}tKUeeC&#uL8 WOy�>�|�5��z�Q��W?��	�r�	�}��Z�T���E����f�0h܍Md!\ܩ�hD�\R���Q�0�ʭmS�s��E3G,��'��;wV��vgk-��)Fp��ZX+���i}ec�Fǃ0R�j�v�&���K�'=;�.ţt��5׿���	\�/Cީ:�kϷ����?�q��c��+��%æ>o	�*���Id�,4jABBõ���Ϗ��,�:U=�M�*����2��:8�3�F'h6!��� �p��m���h�'� L�B2l��lUA�*xd�W�$�T�,�Aߩ�؛��n�БhS%�{)➺j�j����g.-��]� ���7dܴ+Sơ�;M-�ǌY�����2�xp�G���B�qxv5Tt;$}پx���j:�jJl���ޚ=��-=�N�=q���ZཪL+r鑅Dy�j'�Nf�F�%6gAk��u���5q��Yw��G��Ɨ��5�%��mN)��������lw�,���t�5���d\0� qF���5S{�V�bi�Fmq�1=j�L��n�Py�O|���m1)�N���������@n�z��m���u^�����c6YD������3�vm��1~��@�^�f��+>{r�@��]��_����c*:H�1��^ ��,Ć�;ș�gW����֟�ì�U��t����ՓEd��~�e8�:�$+` �ja�C�]�����;�2aM��3Ұ

o����H�Z�ʏ6�\`צ� �e-��'�s�7`����n6�0-T ��̈́��l1-��Z�l39;�ș,:W��� ro��fA��U�Sk\�w���8��@$1W��g��w�`H'v!�^��Xz����Ӭ����*��'�>����5�D�rh�ݥ�!3b7��<B��^(�@w8�R��"��+wڱg���ry�k��0��O�s��K��[�
��)��%^&��'�k�e0�	Q���]���ψj��	��
Ş���"GT����z���c%4�'
Ԓ��xN���?�>,������/���,�CԂ�l�t��#�6<q��� �g��I�D~�}Ϊ��ǣ�rIytB��_x �����{���O��\��rf�e�7ej;��C��)m�FɌ��⍖��2�pH�`b^`$�7A=��q����8u6�߈b�0_�x��#���ufz��`w$9�+t&�����3L�+V^˩��'-�0���vɕ��b��AT����(Xu��}�x�mG���;���
5̪�?j8�6����rHS�����	�_6l�{}b=���F#�d�L��߼��_��?n��p���V �A(N^hu��X�ue���M��P�arW�z��� ��p�?���߮���ɗ=�f�]�ưąj:# 3<긲�����CK�a��:A�V��E������J�ȣOW�E{�%����2�M���������i5��
��c��}�a	O� ��Lp7>Z0��!Y� �{�n��Z[�B�V���~ڗ��\1x��_���M/��Ф��y��W$,R�ƕ8f͇����p0�� ?TV�<�6�J�¥g�h����
{�������]B�N�C��Z�>)�R0'�l ��W����r$�J��Y���Y���j؂����q���'���mB�o��>y��w������3ȣg���`/�9�ΰGk�X�{�>5 ��JT����&�G�(	þ��;˻#:d��Hz�J�"�f���q΂^e���G��+:������N�:���xڔ�&穤U@���
���7��B[����c�P4��6Ӧ�d#��9ہ�[�˙q7��W�u�7]�ũ�J%�4���9o��iz-Y��z��.l�X�_R�)Iʀ����F�����/���A�=��zM0muV��_S+:W3&r�1Z��x�D���^�p��� l;*��ހ�q��f�����p��6��J��X��߉:��l4A׃]irWz)���4Hdv�am�^�t��JJ��7V�� 姦E���]�q�b�pn��u���@v�<�<�f�\��7f�g����AmꟶB�j����P3��W m����������x®H5����){)k~+�YR�}H�t"�����GL��P>P�����x+ۈ��b���1G����f+���VO�R��/j	��}�7��o!���O�ʥ��G���ĵ51��~������#���L7-�3��@��̅�-�[f��H?ޓ�;T�|ak����x���x�ۋ,Ҋx��0��^��σ�v맢�
��۴%E��L��i�-hT�}�Ϸ�nc�i�����s=�2�;k,�1f����K-�u���oz��C2��M7�0X�����S'�*^B2�ĉ&
/g�Ɖ(�Xt�����Q�u�ˮ�ʿ�`���M^H�~��<�_���ߨ`)��S�kx�G�R�q�/J�-(�	�r�����G;���M0���c�27��錺gN�x��~X�����7~	R����N��<�/j�hn�|4����N���`���Gzh��Ư�����4�e<�/j�SWv,;cSX��! ��>�Q/y(�ڹ,��u��d�>AbJ���WI��s����^Pݺi\?�d�L�fT�<�$ce0,�&��x��d��aZvy,�0|��+ǚ���-<#����V��Q.L���bhڈ�v���}���4����V\�����Q?��gFgT��8�m])_}��?M=k�i� �Ob2�xa6��wq1����&�sR��0�\_}Sjxʴ����S��W5�#��^Ƚ�=Q0����UF�JNK�7� �+�vJf�J��
"Of��6'#��gU�探�4�r&F����e�y1h>�Đ�f�?\�s�	a�q�y*��yL�O���wZ >"�|R��;��A	��j�H���q�Iܙ����$�����+�0�5�
���qAc�4����S���Bz
~@��,�L*@z�0�$JZ�E�j,��A���f)H������8��:�k"����'��?�q\S������,�����y��-���k�X���L/N�`MU;+)ґC˪�:� ��!�3j��=�˃�%�ZV�Ԗ�����q����7�>ήl���_��$�!�>����̹����Ș9G�GAs�������t���x�!|<���C�Tme��o����+~t\8h��ٓk#�6�Q��唣*�p�J[裌�1��"< ��3��#,��M����8Sm|�9L���J,#�����g��0��9#���9 "|}ˤ
z<�6|K%�N�g�»�ڭ#����*Ɉ�}�9����,�ţ����\77��(x�򽈕Bjh�1�Q��I�]��%R��5Y?#w�Ϳ�M����י�=�������|��rk)/�zڲ�W���m�i�s��[n��Y�!�w�5��}ǢcZg(�5���_�{�s95
�XJ�g)P����넾l� �36�X���V�X2{n)�	��0D_����k!^����.t���b��$c�Y�#ғb�'��{��=}��g�E����&,2u�r��H�:84�q{�`�_��p��@�V�[C��l@�*s-Y&�i������ì��5s#�E��hTb�;�v��ZA�O�U{-+���Yؽ��e�裖���=�3'V���$!��}���8�9HS��dxQ��ɥF�Ju�cӀp�~�+���T�TDRT�,��4��F`N��.�����↎tP)5 �4����%8�O3���F�*	{��0�)�#��-����gdZ���g:��2wfL-��f�eP68I5T�?Q�;�i��$�X�b"e��eJ�?�2��	�1����s�a��8̭�����%�D�N���9�V4/7$�Gu��تK�wB!��je�d�������,�ԍv�>&�!�P�0Y��q���ר���(#uN����b�����]�U���a\�O�/�!�&ێJ��؎���5eQ8}#��d�}����l�)���s��s����Ų�����b�|Q�F�<�s���,�y/�h�4:�ۖ$��ވ���jC벜r����UHj�)=�P<�g�ya���-UKEL6/��2�􆌇�[���">�lcO�Snkl�Y���&Y+X�ĝ�d�@���^���f����Y�Wذ�vQo�k��� ��l��P<��D{.��s�>匟�����XW�W>&k����"Y��J�	�n�Rϭ{7�A��Qe��A <it�X�F�&�3"Lќ������B���x,�}�2����������|^>=�k0��˓e��Rr�v�Al{s�&��Q�8�P2?DXܴ-�-'����d��c�>&��s���牌�ā���׫ӵ�zC?h�a��N3�Gc����F����|��������٥2�K�-��ߞi��e͋�e�9��%�	���2�؝E�!L<�Y}�(�_ֵ��h���"zq�bPP��*٘��1o~�>y�l��gz��{fj4��j����5�a6�s�Y �3ֳ:��ɕ!��|���f&���.,���Cȿ�^F7b9������KG��8<���Gw�~�� i>�F�^xf&2�L�A6���(d��0��6��L�/U����\�>ʷ���-j�[a�H�!)#%�r��c�=���$�jX�z��X����9ӥ?U����tT��GЗ�1��.�8�Ӌ�� 䝢��CB��Vgru�-n���DTeq�o�����Vgu���V�t ��L�K���M(��n'�iJ�����H������1�D����/jk��A�.�Ԓ��<����[�S����q5PQ���+�^l&]���6���c��i��eL��I��l�R)�[��-J��<)��鸸��n�d��$a��J�ped��0�/"�W������Zϡ��-�bE��C=y�B�kAr8� �3������^+V�1���Fq��N��#�i�Ҷ���W4�a��V�7�~wu�:9���:�I�+�J-��1�J!-R%>FA��U!�jZ_U`�;��`�������N腊�.�ϲ��Bp�,i���{��%�J�XY�mUn}�I�lj���*Ek�WE���r`�f��1��Yl�~�nT$K�V�%0��\ؾ����0X���)U�U��}Q�kL�ܟ�#OQ٪}�yͯp�+�tڎ�,>��Į(1��5��4J���pP���W6Y���d��I!IZ��<�t�\B�0�!M%j�[�͇,���m������{�Ud�]�V붂 uW���JW6���ũ�����I�܃����ܥ8߸$�����^�YCF3�C�AC���xJR6�*��O)qc&rD)G�uo�J^ܸ�"|��Z^d!�.�]Մr)�g��n�{-���Ǽ��M�|�rNԝ���)}�`��_���k�y��!�Q�N>����l���]���v^��M���mǷ{�{�Ѯ�q�3_�w��9�M��~"�2����DCŧ���r*B<�㼵xgc2��i��u���Ԋ��|�n�@�ј�y�Q����Fi�|���޸Mj������)7t�2������M��]ZP�[����x��ϊS2�Q��.�B�FA��c�8�2�e\� �|�+��
�cN���&C���~��\C�c0eL��6�GW���d��@���Qa����x]
�C�.h��Y��᜻.�s��"Ўr�XH��'w	����s��fm��_�$�5�ہ��[:a���pbe��G�g(-ga �pğA��y��j܇���+]o���S�`�a��.��y�Ǟ?��.����v;���M"v!�����ƫ�ٿXB�+3���/�����QS0�PO� ��&R+��{�T^�%C�v	��r�Z�`a:ul��y[�?8�ǂe��jc<8���i~Z'hm�}4�L|Ru�9�b������%7��"D�+�Y�!:S��\ݲ��Q�:��a�	U���o�96Rn�Q.����,w�Ku��,J�S,�����q���&j�-�����d�L���=9��U]��N�;����"��m�Jh��E�*����<�(��^�'�A����N3K��A��{�z?�Y���c���5��r��6�FX���S���U��ǜJ~�6�8J�-ͤz_�S� =kY�	x~�,� ŵ6X�\~�#g����I�2��"��i���?ƥ�����3�B�3�8=_f�
�h�H�3?�P�ԉ�p���Ԟҩ�]�@��c���h���e��������=�t˙��
<��T��w V��#7/�n���Eq�ξ�X�]61�/"�|�E8u��@����;�ސ[���׀��<=��*�N����H2��T�Q�8s{f�γ%;گ�LAʹ��3�u��n9��j.�"�b��XIsse�KD�N*��:DM�Ao�I���WZ�s1�|U�!��Ɵ��枿IҭAG'H�c��SW΋��&s���/�e�����(q���7��)!�zo.�a��`1ʄ$�[��a��H|����Bd"w����u�0������Mϱ�CU#�����OQ�/��`¤'�r�c�[Ƿ�a�����	Lմ[�yk7�M`$яR�Q曧���'�� X�/3U?���I%��m���j��桙��f��Bt����V�f�zK��q��t��3��o{e�g�J��'�6����h�X6�*�}5a3�ky#��!ӂ���X���4O��i���J�vf/��<��@�����@#Ӯ�M��\���IR#omy�ͪ�G��y�6�dO}��D�dW�݊DP�%�!%2�P ��sy���}\M��#E��z��W�5���1��H���Ʀ��S�q��p�B�:D?��9���k�HTl/\UO{+_'����i����C��^h����Y��/��cVHQ�v�kG/��"�1K'.vqb���i4��h|��WHj��>C��R�E����G�X�
y�,���~��@1ԇݜ�;6>���"iФW���+n!C�v�� oy�����%���`�Q¼ɟZd0gj^�.D�ؙ���_0
|�5E������cs&cɓ��UX�^�[���g�� �2�?���f�#��t��*gg.���`^[.�!&�7��U�4�I��8�h�&\_C��q������=A� }m��gTdkʣ($։�o$��X5�����X�(��_io5qL�B_AW넬��R����IY(eXW��|:Uv��Ɓ~��k�,�)�a�=�|���uUC�1�0'��Dw��?��&���$�-_��>��I����������Ņ��_N=�t� �*�Y��-�=��������vl���ؚ��'�cύ�`��)3}�Л	�O�d�C|���_�V}M��ڒʀϸ<���*��^\sOYO:^<�{��՟dصK��;�ظO#����� F�����h�	���ȧ�Q����b���k�Б	�%��t�Lk����M9T�^I4_T�g.��]�[)��%.��0�� ���L���gօ�P	qC f���b��G�<��S|��_%��5�e��ݭ�&�䪑s�:OOםCLWx2�j*�C@Ґ���]��(d3#��IS`���喇��8Հ"Ԁ���������x��k�����?�{x�On�8�'])�7��C:�xܯKp��OB��l��g�`����K��A<�F��D���j��͒���e��u39����̫g(���3�iMP#lj�&�X_���ۀ���JPe��\'��BO������Ը��Q������.Rt�^�w�F�6j�h����e�iu�-z�/��4��͈I��Xe:�O2��V	PX�Q�QȐ!����GLke�Ơ	Ёi�pJ�,>ӳP����8D�e�U4"��#hZD�;a(������	s����!��$��MJ��oj0`�h����ގi�9�
){��=�
�78���Qa�8X��iZ���B�i��O�%�� a�N۴/U�w�����W�a"�~�]���uyȍA�4�`[��|�K'�X�67iHġ���䉄cS�������+# Rc>H��T��}ŏ�u�ȡ0H�Ζ���J��U�T$�w�U�$�Hx1=���爗1�Ȍ�	��7u4L���;�y����w�'�D�!����c�K9��ҷ�*�Xͬ�d�(��nb��m؝h����%�dS|n�RI��{��]��Cm��eQ޽F����A&q�[`
I��y,�e*���r��������	Z� k��TBf�IfJ��oԨ�����ɩboL�����%��Q6^>l`���nN����}>���٭�+"�T3�X= d�/�E�@0�L(����l�$��
��Xa�c����ڭ��,�ܘR�v?���()����@����\����v�8�R�.kh�fS3 ����j�_q����>_u��q��U��Ĵ���B	jppĬ%�9��9��o�	�$ŀ��n�PLm=�Y`g�n�+��]�hr���&�|�z����%�w,� Pd�\����<�mS�I����μ�,��p���9R:�	^�(�����Ѝ��k�6�����]��䒝�{����u�870�9֗�~�o�+�ILHu�Pi����!�:��m�T#h>�P�bmc�X����I����:�\��clݍ��Y�6�:8��iD�#�$�	�)�U�y��i}Ԯ1_M3XZS����>�}�ijm�IÆ��1��E[,t�WZbY1�dF�yOST�2��
�iq��km��{���偗�$-_��knh��`��Z���UW���gA�F�Z�O7�����\ӧ]����u������$1��l���FxPà�0�bW�h^�OnYe���W^㖷�l*�J��ѸΈ#kP$�j�[e�ZyL9��.�FQMJj"y����]���f:r|V}���H�k�7'�"����5[T[�� �u�s��@�b�h�5]#�q}ç��l���;���>^9�� �,wm����V�D�Y�-�-�~��)�&s]_1=Z����"�rU(pԐw�\�kl�
u�K��=X��F�8�ؾs��v��3�8i�����\#���hj����)��G���ۂĵ����	�O'�)���wT�i/o��4�v?0��G\)�j��B?�}��(�R֜|~޶&�*w�Le_nCJ�x
g�˨PB�L�����i�K@�&��y>��kN�"�_�:^�f�tj}eL{-q&�2�} �Bo�!!��5#S]�_��L�����VL��{��巹4�9��MY"�E��߇4�>�m���z�uwe�?�{Xc`�] Da{���b���箟��1��B�S�`�E���HBz��6D�m@(�4l��SL�
��BCk=������h:
pnҡ�^e��w�&<xX��N�gU��qe�s�j2���D"���_-)d� �Fb�s��6��uعjK?�1�1� �.�y�gea����|c`�e�d==�R�i��l��xB}4"���
�`��]��5���fڴ���y3k+ie���f�F�i�}�܁����JBK,����%��p�+x[����vI��s䲐�9hɁ�{Xw�A_?}F��t�9S��[烍b���/Fc�L��s�.-;� ��
��������zC.3��:��#�/����7��A:�d!�U;�&aBi.�Y_�� |J�:G�6cO����Xet��%4l.�M����rb����M�dt}B6r��iӶP̭�:�.ު�o�am�;������"u>*Z{��K���Fk��J���<�_����;%�"�U|�k�N	�q��"�=�]{�̝��1vP��tkj��	1�n]���4<�y�i4���mr���e?U���,^��r��a�05��j�{Λ'��~��j[[�1�1tв��Z�	�^t�����W*�ь����B�v����"%_zV�-u�����WL�,�W�;��[�L�&{p�"��`N7�Nb}M�).5���SS���l*f>b��5� K��H�`k\1�o^������WϮyG��� ��Cg}�خ_Ǥ�Uv˘�k1�vL�Q�P�ٍ�1Pi�S��va��uM�����=��׀+S)&��Pt����w�����yk�H��Ћ��A��cogw�V�dN͏�O.��d/�b�~��k�T�l��g�e��U?�@�� 󾄮O홑_��˪�o�O�%��}�T�u�
T� 4XڀY�>��]�uM���g/���_+���BAI��q:��.8@d����%�a!�����'d"[�Z�T�� ���ME=�iy#����B��iۑ�ǹ��t�a�Qj8�w�����橩��()�Lu��r��ڝ�]��a���<���Hǲě[�y�7K��@16����n.��
ǯ�A֜	T���{4Vv��	S�gM�"�k'�v�黳�W�a�ߛ�u���t<��i���,hĤg$rp�ԧ�$AH8;[K���P��Wf�Dn������X_`f�g���J{𜥊/���e�ʊܭ%2�bPq�e�.�y=��(����! ��n�f}�Bg,Sg��sP5���=1 D���9N��ʁX;�S���M?$0wvX��Шz��a�l}e&���
��!�����kr�.�N���{��,�s�~�>��m�|��s4Ez��4��%�>�/OEQ�/Ax5�>��ӯ�o!���Y_y����oU6X-�\����Hd`��T��ŝo���2��b%�`9���3�ͷ��:@�t�|oIBU���+��^_�Os��Ŗ�-B����-+mo=���dN���˹��J�ތ�4��3��B`)F,����Z\��O �^��L�C2�aF�� �"͐x�[�uJ�kfu��@ ?�lB��Ĕs�M�q�Zn`=B�8|+�iEp��mb֙dtP���PkoP�d���w�T��9t ��i�����
�׭������������s"s��fDiPp|o�y����?n	�,T�}��y�*�����k[��l��W�d\"��qD�k��s���P�6K��B7�L=O�.�]gOiL^�J�n���D�gZȷf9&xE{�E��E���%��,3��<#*�}x)8�@A����§n �z�F������� ~��3�>�*A���Q@Q�_?����߲+\��H�Ć#w�Q6�I˼M��;�P�>(����z��yl��n	���|%���?ƔH,e3i�~�*�-K�&+�F��n�A�K��)C���žWdfg ��6�����t�VD 4zx��ز#�F�k��]�&�7�|U�y�cxe�4�(��0)Π�m��	��������nD@H��9J��?; �W��7 PbkI��4m��lE3�WX~=	��ïh��d��	A�2���K�y��x����#����ծ�E';'��! [�ZV	�㲈?���@��:b�v��)U%���钵h-���ӫJI�gt��bc o��~�[�)&	�La��k�� Ԇ�f3�O9
�
+9#kiHAP�u{B�'�":Bs�r��0n ����������� ]صI<�<�wQ����������*����S��#p�#�R���q���(v��ID8ІZoz�����~@k��h��SUD,�IjWZ'��	���А�W`��liwL(J`I�:�L�k��盯�ƫ�W��4{;d���k�Us�xa�~����Ĉ���V�}@�TY�j�� �1��=��(6a��.�O��	P�H
«�ys�n��x2����X[�Fc��.S���p2�-�	�i��g�����n�E!��T�Y#�i����#7خ��=����4���v�� M�l}�M���3� ��N�>,.�:�G+_�Eg׷K ���x������ Zl��F����=�F���R�l ��V��u�6jaJ���o�;���)���t�"X�fՐ O��K�?]�����cG`j��bSO}ߕW�.���G��Ń����
P�2�������by	�ި�7!f�-�	����5F�|]s ��?�����x����[�Ol���(�����I���Al'��ђ�R����������N��3�r��4m�A%����r>�����$>>��l>�co�P�)hJ~���U\����J6d�e�)i�?P��$��76mQ�3�"S�)�	�YyT���cW��E	h�x��8��c��U� ;�e�ί���@�]��ѓ�"K&U1��n�	�N��}�)��ng�U#��}�٘@��=zsNI��m�¯Q��+��`u./�݈�&Q
���bϏ�7XV4E�o_a��8x��� i���:���໚@Zn���Jܻ�t�O3�B*Q���HC�$�w��>VVa���I����o�9�1E�"��\��1��V����K_kY�Ϯ�PL����Wy9�	�;�g�}��b�fYE���n�<�"��¸[z��_$,�Aeϸ���h�A��zG�9T�H�
�\�X��;����Q&�#����RF���B�ľE��g�#���i&���ET9�̃'�W�΍�	w��.�(��Ym8Jy
l�I�^���ʪtz����)��N;�^�����D�YO��H��7:��I������{�F�?ԧ}��*Of�L����ͪJ��٘R&��B���O� ���t{|�B%aV�ʻ�]��I���xW�n�h�镞�>�}�nH��-ZŷU�#�߅L0��@aV�.�3~��G&5 NRse��D�)��X@j��/Rч~�ب&Ϥ��:�z�ޔ�y\:����'E靧�\Rh���)7��I��e
e��c���꠲�2�W�L���2�o��U��Z�K��O�Rk�����({�W��hH�M.��R^X�~� +(���ϗ�E�ml�VԌZh�;̥�%��l����
�C=���.KQ���M��ݖ�6m��P0��J>�����xG l�&��,Y���7�?�_0W�.oM��ߩE�V}����p"#���2�@��e�� &=(�bO�w��@�f�Y_ZD�ؖ��eIN+�YK�d�H�nW�}ڊ��*B!%K%%�U��P�!K�&������||��'54�2��j�<?�����-;�q��r��9�����"�IbJ�j$I����F_4X�Αɯ~�V3�� PMy�������~�����/���Qs���2� >�t4i�h d�n�30(��Ҙ^AuҀ��U'\�i�d6��/{R�m:\�X]�Ha������!e��fG4np�P�L(��Dn����Ƅ6k L���W(��3o߃~�ѥ�矞Ws�s~?���/5's��-`\]t��;UM�+�2�@'d����]�X��q�f����b���_��:����ĸ�ן�l�}���P6_�5Xʢ=.-ю!��­�M:[ۣ^��3��w��ie\0�$~$��|sfR|:E�_&�<�p�Ih������E��$>��`szP�/4�1�j�-ͧ��Y� �)���Q�jC߹ԁXx3���1D�*$�+	8!^�N]��:�]Fy1�BD�$�*�[�Q�
�Ru�q≎�Χh�+��U��Y��Mwu�����ӓ�4�V��b�"y�ϕ�����F8a�w0U�MC�`��6I[��
0�Xί�!w�THe��{kf��%�2����i)�~j�~d�l���v)�$�P��%��2��<�����U���VA��Ӂ\i�n�$$�����6̃�jB�{���P��Eo�b�¢��l?jmL?O�(w���@PBa
GOY���8��±�k�Kn,<��R���[:�+|9��R�0[�qw�%�|D��n�J'�=px2�n��}dG�đ�a�ȶ�?	FN`}-9Wv��|~���9����aE���a�}tu~�kt=D��2�(MbvY-��%���O ���*Ea��O�/��^�#6���L"�Q���>0�/
\}dfkTK����|����U��ʐc���6���
�|" �@�#73������6|*���[�K��.���vv;�2n��@m���v9��F��tċD�D\#=��C�v�ڽ��j��֜�jK�rW�I 40K������'��|��Ѿ6�=Ggj���+>?���#��
h��`���r�f���}f�Ȱ�j&Ffn��A��M�� ����6}X�K��op���
�����جj%������z�e��k����$)5��4�k�-u�Ȧ�/�҂ OFQ���V=���r�]1��w�rk $S<]&��Z���#�rc`�� &������q�y9�~7�jy�B��UA6>:�-�*�Ÿ�A�Aw���`�32��@���?텸D@�fo��4.�d�MZt
�+�V�pX�N8j�œ�?E(�s��2S)DA�/��K��W{K>P��R�w�*�]8�؍���;�2s��($��([�j�5��]�h1�'���M\�5@!�v'�J���ëhaF�Wd��M]-^������FĦC+�Ҿ'�7�5OQȨ�zw*Wc_�gȯ޲	�x�So|�ih��X��q�H��9x�H؅g��A���7I3�Nvkdm�)�쓀�t@;����R�e~4��O��`�r�~�VD&v 3(n�7�n��U�"��?1#�	�k����A�֘'���/OA|���\�&�'���#�$߶�A�a9y�LWH��y�n��vBmF��!�ٺ�����(F���HͣC�)g�w%b��n�O~D�0�Z4 ���0�*�@�U�|�\�בT��d�{�F�?D����O$�{�!}�������sƍqΥ�q���5wcI��3=/�3�����7�;"�Z�����㝞��]�`i��J�O��w���O�a�U}��.��)�znNA����A$�)
y�+��T�������]���4Y���H۬�ǝ�i�s�n�٠�Lp��Sڹ_��nl�ؼ'	`ӶV6�����T"�s�[/s^ �#�A�2�{���g6��'��1� ΁�vv�<m�������w��bKJ�+�"�6�m
���ONV��ou����\TxCSKޮ��^��V����/��N��Z�?��K�}e�8�:����zGٸ��ue�M��폚�B�e��\���;�nQ�:pԻ�a%������`��d���>	%��'�-�Tnj������'��B��*����Ʊ#�JQ*�js��,�X ����t�I�'E�[� }�+��;�ɢ�?$xXh��Xڗ��,�	���B�W�0����~GS��ةQ�J^f�
��c�.�0������� ��J/�C�OP�+X`@V��5@�sΌ@�0ߝ��2HB��,�ϊ��������5�3X_%_SK2_cS>�#�X�]�*���t���S�|TI�`��&��ȷ��M!CP�f���;���D�^�%�:�f��
*��ᄃriš�f��1#8x�; �Uu���Pc@�?U�W��\��.sk=��&�F.����p�N`�(Q�-�Vu�ٺI׾�u�A�S������X�G�[���!6a�����Sa�\
�m2��vw��S#���a(��C'vgCdc��"?�-�M�!r�ѷt�uWދ�݊��G��2v�������#�4��7�<Z�2�oW�{���Aa!�*Z���e6E�{)ۈjz�)�/�
�(3��"?*_ʸ��ʙ�?��K��1�3��yP�7O�O�&�;�_%���JלV�  }��褔㘱$�K�&
¹����;�c�J�zr4�9��0bw�bē�V!d�죎c7��1�,�ޞ�ts��
eY1��r2���$K���5b_��Ȕ��^�G��v�
ڶ�勎�,4R:������G=�qC��J#��~����g�طP������A��a�
�җd
dڝ��Wٚ�=R3l��z���پI�wA/��Y�����޹͈K�M�T�b��Rk��F���D���H�#��8��MF�v~�'6�MW}j�f�Iv�Vho>D
��B�o�zQ�v{^|$�(|�,���0nIŪr��HUV{��줨w��VI	�>�"��(���۹�yu.�VD�j�.�d�:��vq��lvڱ�5�)Տ2D�_Pf��R�;J�F˳�A�?x�űz�"@��y��w�q����N����!VMe�&�Q3�#��H��A^��;� ��v�_�ԚH
S4�����r ������6N�%N�%�j��T�+J�0oP�e���_�w�WM]^���2��)�X,�p�E�ؓ,	� �(-��Vʍ�Z�\o�P��}����K_�Zp[X��S�����Y\�����C ��tv��1,�����iq�J ћE7V��ߩ���K<��V�أ0�m�ս�ɑv�[æ��rN���fk��L|3p$��)9�U�WD�{���(��_���f�b�`!W������zv�B�����Za��N�T� M�H�M\�[�T�X��x�c�o%�|����fQz�D3�Z���K�`_~;Q4M���8���̓��͂�����(�&�(6�,�B+��1���*����d'ax�3���0���ISj�c֪��G�c��e)���26�"�+�W����"�E��W\� :���uڍi�LX�_0�s62<��S�\�8��x�(�h �����)]�<,��r�R���O�`F��hU�ж}���r{."��5Wi�:�Z��8І�������JӍ=��d�Џ��KnBABW��ăe8��z>z̨������sX�F�e/U��ɯM!UYiu�92tw���۔.m�Nw@���	 is�`�tq�
<�-l͜��\ӭ�'��K�+���a�dtox���(�5��9�-��u+�_s+p>y�1�.B�N�	�(��<�Fޯ����z�?���z��vR��[�oqi� �����[A�y(���!�i�+��D�Ұ�M����/�32 =�*I����ڿ�A�%�_L/�b�`WBݣ�|9��~+i���`�
�@@S�īb�������e�{�]��
��'��n4��uq�@��3�ǯ�{���
:���i�m��G�^8���F"NCX���d�Re��)����\7�V��Y�腥&��Mݠ�-�[�Y~��ݰ_���B���uI�ꬵ�Qg��:��7X�u;�2��XYN��"�5n�n������Ì�£���Z�{�oW/��}�ے�
ܓ0��c���Ʌ�\�8f9ǌ;�q9�"E�Eat���|�(v�#<T���9Ի$4(�^s��Q2�m�Bix�(\���
Ĭ@|{�QevD4/SS��2�^��8�M\��g)Z��O��8P�^���Ƭ�a.������9=�Y�*��̱ʁ3�ax�=��)���@��Jh]��:��>�)rjT����O)8�E�y�}��3.�;%�Xmb�_�{DW��W E��vwh�zgM� ��y�#���>�ɦ�I�T�ς	���t�I�Ӯr�k��[�>�c�W��������Z�ӈ���p.�c��]MRѩ:��796�$]_]�4o37��0���G�d��i�ј�!��:gķr`�b�Cl�[�b�Yd�}��}l�;h$X�~t,ݎ6rHoyI՞���'����u�l�����1���eG�D�w�lY�1��$�L��լ pA���E�2�*��p5�`����3,l*��A�4F9��U{^��.�Ic9 3I#9���g���{E��m�KQv�/�
�P�X���1�[6JxI=���c���gO4�~�]�zx��h��Ȏ���;�s������ K-���:�:7䑭<����C��҅��a8BmxG�nfzH���T+�x#�䂞j�T4r8�*(���~~q���?LMf��n^��>^���(�1���j�SF]�Ɨ��u��x�$,���hNrmE�ֲ��i���<9v� ��c6e}h�M���f�
f�(Qި�5��˽[�۷��a����z����T�p���Tۡ��������n\��`��R���>M�dB0R��*�a ����\��o�5��!�� ��M4�'Ur�����g�(f�w�6=F�_Ax�4t��r�6L��� �{�pϡkw�{W�¶�A��@nu8��S` ���zǃD��*�Pf��b����z��?��u��_Nx5=Z�Qƫ����$NH��{~G�Р,l�L�>�F�%˺XI�_�ܫ�)F|�W�ǑIJ>?&��e��7w��whS��:o�%�ET�3�k��ǅz��"�b�߫,�h����I()��s�U�x%��ܸ��눾 ���1��`�3����e�0+߈�����������eSB[�)�n�*U�,�O��Z�v�kv'Ƙ�~j���n�?ܡ��Y� ��?��Jd 7\~RDQOP cjR�,�f���ͷ47��.��R��j�]}��7���r�/���$ѪN8Md�B	x��mΡm���v1J��k4M{j�^�;��Y��U��֊:�����<�=��bn�]�#��YK�Zv�2���p�ұ~��B�ؘ?�D�t�va�c�B�#�}1����ssݪ��Y��>0��L�jLWEG[����r�7u�8p%ݝL��������`��|V	#|�on
|&UՋ��di��i�Z�ݓ�
c ^r���m�7������0�-�R�|�*��՘ɭ���p����v�D�)����YOH��.§�����V�W��ʢ������,����X�|o��\f������9�D���nfl�8I[Db_,�3Dԝ�RE�J*4>��g;���AW�4�b��0���_6����OYo���0�8��U)\p�;�a��D����b�����U�o�"Q�3��c6;����wwEw�!��ʞ���q��m`~Dpm|4���OE����q�$V�M��������:�������Kv�[KV�.�iK
��:8"@�cR"XT̪�\Fd�ݍ\Z�g_UE��RGBc\�t|l��h��b��X�]j싽`�N䇢K���>"�;������#}v�a�9^�|���?�ڛVN�
�����@5�A;ҩ���#��]���:����
�Sj/�0PRQ~�cy]�i��ۉ�Xz<�8��Z���)�B[yGG-�.0��<*ټĈ��5"oy�n�����<�I�gUI�'��W�Ϗv����Pf�/
ԡ��A0�z���C�݉WװSJ*��t�����~:�c�j��F?&�!��G��q���ԙ� �AJA8m�}5���B�?�^�^¾������~���'�C�U��*�h�~�����9��	��ˮ8pi��ɐvS���ĆE?�7l�����y<�䰕<g��F?��\fO���6V�^gN���͟V���D�B�L��L*�vy��w6>��j"D�LF6i����n�ujg�G@� ���p�m������f�!#��P�2�ZE����sW����Yu�kyF����h�U4E�A�L��%�qF�����3f-n������h)����?m� �
�9���A^�2�Uv7r�:~W��-q3RԚ_~a(�r�K�6@|�gB�d�Ip��nN�n�)/�-�S�~������0������2��Q��ϙ}qv7�~+%�pt�9�R��O�|s]�J���Q0"�]!��aD4[�{Å�L>��Y/���U�|���d_cU��*�������|xF��Pr"Qp�/.���'�|It#7X�	���^-W�Nɜ��[�H��J}�9HZL-�1>R7$�O\F��Df�B"��G��с^�j��9P�;�
ס!i�kN��K~dKc\�W���	���1@\�A��=�7��$"j��R�1�!�/�@d���Щh4T�>��#�4t����k��䰮�3�@-��gֹ��d��o���J��})s`��)������iȠ���ө����x�K��Cc����+%�E��xĊi���0h^�$�^--4�\bJ;�� �*�$�)��� ���FZ^�����8/�r��Cf�64.�����n��c�Ɉ��p̗�9�|�]�_�UzE�Z��AHR��
�?���������rp�]���O����ʎCw�H�̉�(q�VG����d�RD�ɕ~�R�J�@���� ��ɤ����[fv|�4�E���Mb����]��xV�b��P�y������iTT%%?�[�sU�'݂����=�Ađiծ�eyȻ.�B3��� �.˹�MB=��>��K (a�b�<G����� ���^��dc�HP�Gɿ���9�.q�B7��*:��Nf�sW�x')�Io���Z�������f�5�#����0\��U8�轲�I&�;<+nP���CN�Qqja�liD+嶛�X'��8��� d�[�%�����3�,����V%�7_���֓K��$�̑9ܬ-�YK�R�_���8�~�Rq�;��z���))�(�X0I� ���HQl��#��۠�z\��Π��/4�~-~�b��TTn��0'7����;�ڐa�~{X��⢙�8R�2bm=\�qH���+5��M��S��3�䧏ROr��Yw��je~��yeC��3�>vr���W�GjM�t�.| �d����P��Q̡O��e�*U7�G�*�=���*�>\�����:ԡ����XY^&�{l��PSd�R�9�J!�`���-��O���$�,�3��4��Q�v�xs�+�qZ�e�Ag�/F�M��-�����m~U00�t�s���UPѳ+(iĔ�6D�q?K��h�hI��`��.���#d�sg�_�m��<!I=�����B��FML?[j�!�)K�������C�����aТ!��0qi�q�����������c��ܢ�$\F?���E�~��<֠@�]K��k����A��F+�L�{�w�;��[����
|��xG�t׼S%(���������?�4�V3�����h�EgR �>Kԩ�^ǎ���b��Z^e�.%�"�v=o�ҀɅ���X����^3څz��p.���M�j�JDj�6��C(�q{�;��fH��o
W� ��厔l-_��ԅE���o��HmÎ��5U��v�����j�����9y�w��n�'Ww:=FP%�k�`��շ-�E�*Ҭ���Ճ̈́pvx.�6&��Z
��h��r��ބrO�����J.�����=vw�n�G�rt��� _��,�=�S�B�(<��ĕF�*A�����V����j�EM���}�V����''g�j�ބ����?�h�8a������ˎ6��,�,S�*���\j��Z˜V\o��秏w14G��'���^��'"[+8����}�]I K�q"�S<߹jۉd.I��v��9{E���E$IA��3҇\�S%"�L�B@�����8J�AG�\��C��8�i>�AGX��F'��1SДL��<Y�9��t����"��*;��Lh�E/�6�-���;M���ٰ�G�[�u�"�-��pGO����s��\�jBi�������$~�9ܯa\��� +��G�WL����a��[�h��Q�_±7܏����$��\�\�Fk蘋Pn-���޴�Ͽ�����+�m��'s�A�>뽢�M4E2`�Y�Ec�wR��t���_����{x���V�=5��]^m�r��.�H{sH~�f��
&�y��! 8Vr�?�M��uI�r<S��m������(�h�F0�bI�:Qa��Z�2m����xch4��h���U�D����8ܚ'��@9s![��Qb�?���F�uZV~�@���:��A��*A�H���y򔧆oO��_��ߪ��"�� M۩���;�C�b��t�3�r��4Ov��2prK��N���<����ΰck�M%oŉ2�u4�<�p*��c�O=�.��4b���0��E�!��닌yf���m���X=Q�FQ#\������̖ߧL��D)M��c�S��]����&�����2�~ᫍ�����L�W�G\`G��K��s�'!?�j�81��	)+@�6��n{�ԩ�V�Z���JStD�+\'QT��P��a��e��������<c��|�jM����Ŋ��{�� ���i���V�D��P���"J�K���$�9�$�{2k���;"����AL�X~���0�8�,�� ��=|j����ó�ml�i��K����#2���J&��{Yȩ�aZ �O��!�=3�,�7� �)���:14��rmz�=�V�j+�����A�P��G�S|\F� �F f�<��9�Af��ғa�W����*v�����g��Eu�iTnL�3��~YG�  Ta+C�ٻ��3݋�HTh���3��p�����a�� �L��JCj���L�w�'"������n��4{x�.��>�Lh#�R_����=cM��ǒ{0�~�k[�\��S�? �t='�j��Yv�LY��T1Jy��wd���f-�m0A�	9�K ��L����x�BP,}ۛ�F��J6m�Mxm�!k�Σ�說~�O�1o�<"�MV�n�W9��]-=ϏS���[����d�S��VEiH'�>*�.R�/�۱�0L��e���J&����~Z�K��TG��^?N�*](�X6LS�_&,�����q��2]�q�d�p��	���~5�S(�-3lP��T!�/��R�=����.����pm:��y�9׌uQ(�}�I�-�R��Z�k�͑�Gx+�+�����0i�����ɺg��ΏR���B��^����'<0��o3�w�:�0y�Ci��lu�zA�̜���w4���T.xgXIm姀��I�XgqQ���GƓ�ֱ��}�%���I�����$�1l�?<< P���3�x؝��V�5���*!)Kt��X!J#���Ws.��� :V�/%η� �<=#��߷@�&�u�����j�j�Z:'�[PX؝���焾3��is��û��ň�$�*͓w{y,5:�K��z?/��n՟X�Һƿ3*��H-���Q����P��T�͋��|'��}O��Pj �
3k�㓿J��9?������sj]�ƶ\8�I};�T�����ߏ��dn�U���M� ���R��
�|xl,���PZ��(Y��E%I��M_�Ur�f���|P).�6�PS>�� A�����׫�=�Cr!q�A�i��l����si$e8�+�C(��w��s-�/D�}u͛0P0:O(�Yi��/��#�7��h�KUGL�l]>�����N�����G�?�n���<sA�j�����=�K7���Ls�
��5~�A�PH����w �9��f��
�F	���h>�.g� o_�9#�̟-b��O�VD9 {��^�C�F���W]�j�پ-S�;��9b��x�G�ee^^ �d�z8g�QHh��������vcJ���Yb���Iݷ�˧�i�<���	+���\/�m6��Q#m*�6	u0�$0��qg vM	��W���
�J,g��u��2Y��B���~�4W�}��S�lc�TO���	�	��3�R�?^�Q�y[X ��pD�Ԍ�,�-���+Jkڰ�k6Q �U[�Z�?tQ���Tp�.F����ƛ��rʳ���q �xG��`{��������Ç*���l�D��n���|��YD&Mp��>�����m��hHXṐ�.�9<������mK�4�Ddp�9u���9�|^ͭ�J��L�ډ��O�D��J�Q������.F�]�0�L���w�L(���˵�˱�����d�5cyQg��UG9�i�p��{ѽ���@��a_ƍƩ����qʪ�pˆ����[��F[��5U�;����u�=:hY�Z��/����B�h��	��"�8])�н?<����Z�|����%rk )�H��5�ʂ#�2�+�������yQ�u�"��M �� �}Jb�����:���wYLda��ZZc��^-�������E�}O�-�
�g~���虸��͎8)_heQ��kׯ~/���O����a<�)��j�(b+����L
��U�HQ����z?	�H�L�!w��)�%�}/%9�'V�M�MAHz�c�����:���.fb$��S�&�<#T�Y�A��$��M����x�W�M7s���#l�m�s��pܑ��Y�1ћ�^k��Ъ�.�נ#���r8���L��Q�˖��?�L(	YXiS6� �K��x�S�̰�xk���Y��CB%!�I�Cc��+c�t�ɕ�Kx� 3�K|Լ��nO�п>�UrvHM�h[˹F�29�CF5���>/e'�1�4�H3�wp숤ω��fB��+Do)��_F�����?ũQ��9���ւAޅi6~�Q��F�|�O�^�hi�5����\���A���=������Y��>�I�i�'몭��=��� b����J�p�����OZs��݉>�k���a*��j�;oBfR �2����"�(�6i�i_YiOo���O�_������Q��h���'r3���O�Lq姈 ��)���"�������m��%���F#V�Y�i�IH������7@���dG�|�����;%��
 ��[W�UbƗ�ʣ+�8g��X���s�~��O�x���Hl>ފ�3���n:^G��5Y&���VgE��.�0$�@�9	o��㠪[&�5j:ŀd������"Q��m�g�Y*~#��T�d��scM�S:��`��fX�]N������q�jÛ�(�d4d�ܬj<�MA�Q����W6�t�E�_��T�s�^c��c�)ľ�9i:E��;����-����CM�������<oꄢP�u���4(��ޟ،�ɺ-�;�D2y��}rGU��SO�g�+A�%!ᱟd)�i �i'�T�A4T'~��#j��o���C|la2k�o���_�c*%ŏz	��5���]��n#�"[�����G�x�YAE� ֹ�u�fSdB��ɝ�)j)5��m�%�u��3X��T�w,��H���d��x�C�X�|8��d�����`D~�Ѯ�l��ե��29.����V̺`ɴw������2xH�#���7q� �{��]a-P�{!A���u�a��F��D���*#��1g#���0�qj�%�lz�s��s��ٽ�(����r�C�_����k�]�c<5_���#��Nef��%T�,W҃{U�?^h����xs��j����G�?��F}�Oj��O�Y�� ��\"��Δ�Q��s��iS%�O+�C�X��� {��W*���uu�U $T �vţ4�rGF��q�چ�0hP�_A0p�3��I�N��@�>��9%��\�6.QraLc�|f�^~J�� �R��z4��ׇ�d2G��l\�;Aǌ���]8� �@�+�}�C�S_�QsVz����ʎR�}D��Q�L�[P�s-y�q�N��6ڲ_d�Ͼ�CR�cִf�{�}����}�g>2=W�:���z7�9�s� ;@����櫹챦>���H�W���S��x�3� a�����Xc�X4���Y����?�
��8�����6�.Ãz�m��ryH��A�I�������M���'����Q)�/�����!�-Q��)j��Q�_��K=�P��V�>3�jV	�7����HㇲJ���l����U��[�d���{��x;���H���TM���)��oW�0�$F�!�(��	ݯ՘7��)��Gߗ�ri��{e�[���yՋ��)�J\����J0`�Ԇ�������qc LZ7؅��9(\���WWΈ4ާH�1v���la4��u�7>~�f�]φ�?Z��&C*i���~説� m������E�h9#����pa܋S}&}.�����ҽFT�-�lE�E&�2�M�n�Z�'z�:m�X���;�#),��oS�?\@���Ym�_���]F���8�m� -��Qv���d��^���[)1LZOcL�Λ/g��O�H�ª�p>��35L���7XlX&��j�%�|�5G�s�ӌz~Bi6��p�|؆�¹	�h�G9\�n��|�]՞���w�4�Y�@�:�ո6����}jߥg�YU�����A+f�G�6��=\�m9�<����*��sXv{Xn��� !`,�B�]!ND��.�z5�Bd�6l4���C��l�G{�� ��V&g}�pA��;��]F2�'�]�,p�p�fJ8�ڐ}�E�����v܀6I�$�,T,�D:�n���6�chD��g��j����mJB#t�P�,��r,���>Z�z��˿a�����JBN��@�~KZ.���� �שv�r5�hԨ���M��W�����W��é�:��f�&���&e��Q���wv�җ��تP�	S��a��F\�.����~��ŏć�f�|[ �	�*xDn��Yv�����sn"����8eb�73򪣥�(N���Hd8���,�̼$��q3��a�To�ң7�k�2
_�4~fYy?$�r6�CbT@��ִ�Jpے�!�\�ŖO��[��6���I��F���Iv�r'HQ�j�v�eǻ��
��� ��{7�t�g�$Nmϓ����'�w7I�<��Wv]nme��戹�:1�D���E~�΄!8�em{x�,�v����S�����(����	��eЖ�n��.�U��3�r�{㐜���P����N��y( ��0��j��4y9}���M8P%��ek��m��U��ʍ/� �?5]��e1�~+�l=ʏ��wQ]�٪<+�3)`���T;����@cyG�l<��S�͘$��|骝�r�-B2�?b+��V����=c�?ş�[-�b(�+�V��V:��@gT�B5ںde�����UԂ�*lj�t��ȸ��)�'mYjb���ѭT����u�ԋI)}��7�+�W.�4VB�kW(��⥓���#����on2��Y^�N���S�PI���%�N�@���L9U-�XyNV`����5��$:�#7�����XC���n��:�Ⱥ�&�@�I��GS�B�>˔���?��j�ν�z�X^舳��5z��Q���!;��$!�;�Kh��ަ�m4m�#��.gٜ�p��r��27i7]�0J�S� f�p��Ď0T�
��2��\F������4"I�,�n����*:-0
	�� ��#���@���,���<�[U���w�氏��%�o՚���&���4�؏�7�����CZ���#�e(to?1^QWI�F����&@��.�l�l��I�.jm��9;y�m�?�B�)JA���/L�y�-�R�������v9&�-��_1][z�c5sP:�5�'�:�W���\���W[�a��F5�=XႮ�'�	H�FʝTc3�r�#��&�{��j�Gj�D`���{j{����'���,̈́T��e˕(�P�k���Z�#&�;�"6h.Z�'��Ǭr����lŀ��!*OJ��ə�H�~ķ�j���ō#�O,M�o����� ���������g��vh��8��N�B��$�2U�G��l>�30�Y'{n<ġ�yG�o(�\�+;1���t�����LP��Eh�=������U��c��n��5����va��|?�7��ɖ��z���y#3n�D72�����!1��1��2�^�M�3��j�1`A�FԜ��њ�2�ZYM?�Ő�wC�1׊��z�y��I��s�#��C�c��ؗ{nj_�3\%ZboR<���H���b�`��{�T�0�6�}�ǃ���&�s�����k��>�~X��jh��>�^��������������*��1���,N`m�?��9�<�E�,1 "}4{��_j�Ί��p�� ��Ӆk�L��ڷ�}�Hy�yH�T���5:vM���n��o�(�j����ɿ@�}P�)�^=�Q�G�d���,M�y�	,��������8_�mIC�Z�`=;�لd.��l��~� ��(6:�11��9�k�:҄�/W�	;n�eb2J�,` ���(��:w(]����vēk���[��{�B���� ON����e7�I�8��*]�#G��u�]�g�C/0���"�9�W}�8ȩ-~d���(?�iM6�j�T��09�����Z{�W[���V��NU�p%؀O��s�OȆmH+�AZ�9�aM{�|�=PE����|KF�"
���E�{���)��,����G��)&%���!�S�>o��mH�ql�?a5׃EMl	^���%ˉ�-e��/8?�/4����p�a��б!�Ÿ�z��*�dۃo,4>F2���.J�� 2f�*q����ʕ���@���1�����D�\>�YTD4v�CL��9zr�c�x^��0^2t�3��h4�pm�b�2�\5�tQ���;k<�w�ɏ2~�%���;�^���޷C@>��)v������e�W��ʢƮ>1��𳾘}}�>gx�=� ����3k�{���)�̍�_��0����H�I�D�y�ՕU��NJ��6�9�u>��U$��2xWo�~���@,�!��G�[_�6�s榤=��1_=7�9�W:|&�	���:�x��:IV2]�.?ˬ��l��c�)7�c���1�@��1�R���%��F���:=�3� ���B: �{�-��j`�a43`��3���Ɔ��"ц@��ɮ�=SI^� ��yIb�\��S���(�83;��	%��X�B�]U`���U<��C3����|��jml�m�c%���ނؾ��@~�l
'E.T�RI�O4B��d��A�N<-㷤:�&Y�P������zبP_L8|��*GDG�3)������)T��G���t���%�u���~��_x5�s(�g`���J���1�8N;�6 
���Ig���P�<��A3	Z˪�D�D�}�?qR7�q����(.��N�S��?`���Ҷ<�K����K�~>���h�I�����C&)p�b�xB~L=�;_&�D�V��,mT<�U�#nK\�uӖ�A�Yx��l|8Y�D }Y�_��X����)U�Z��c9GxM���-��(t�z9�N�c���m��L��,;A(��߮S{�̂����Y�F����Q4���z�熬�@'��V�w\_�����2���y��:nO��I46@�Gs�.CKM�:]	3V�q��é�ʣ|��s[8�l���&�Os��K���ٛ�ϲ�
gݛ��|���%���p�%&�t��֎�p�"�W�]^�cu��g��x2xwu&\I��8�%+$	m�vҀ����n֕�M�X���/g��z���5��ru��<�`�\����}ju���Ѝ���b��N

��������_[a��w����)�5n#E�3�i�(Y������pC�)Z�����<v|�����7��� ԞJy�K��8e#������~���{:]�{d�P���qJѳ\���1�[Q ��a��ȝ$(�vLi�S�#�/�,�X���+�s=&�:{nw����~M
k�y$�����ĕ xd��ﾕl`�<�1 ��� [=3i���]x�`ʼSܫ5�_J&]Xg����F�ʂm��*���EC�@� �9Y}K�'��|���\�Y5WYdlR�/�)vP��6W}&aV�C��	]}�p�*`0ĉs���{x�ӯx�#O�9ӛ�����kv��8����
XL�P��ͽ����G)�ԅ2�I"*�`R�A#2o���ڏ� ��ˣ�kL�PG~ӷe�m��7�Z�Y�`Rx뒄�)�mj�:.Q��� ������P���-�*:G)�	��$*���+F}�������ǀ�	����'i��R�?�")�e� ゟ�	��R��;2�ܖae+�h$#�L~�w��&	�Nx�y�Jk��L��Syȱ�r���9���&$�C�(fJ[P�H��R*Vv��N��؝Ď\�P~Y�m�
{�݃�|�����9�Z� ���*_�j@��E��7��D��+�e����Y]0�~����:.�@h��|�w����7�d�2u<�x��?f^���g9�;A]�m2^��F}"��j�i��(4��&&3M`F����#|�b���>5E3��ץ�Q�dM~�~ei��A~�Sܱ�3~���?R�̪w�O�l�5p?D�|�N��IĂ��L��C�*)�S
��i��{�H����LX�F��fy t�57�c"m㔰��{;�{�$0���-�jk)ꈏ���U%�~�k���';��s$�����$>t�	����:x@�n�P��`���x�t�Q�9^5VNT(!�gJ�6A*V���h琼㨰�;ʆ%�c���dʸ��4�S�*�`;�:��n�����"Հڥ���'*W ��w�a<������M��=Z@���MiC����� kz����{�X�I�rlHR) �
R���.�y}�����ꭡU�ϒɱ����Z�-]yY?	��۱3��2Tr�?�2otshZgJ%�5O�P��eu�o�/j�Af�Ju�|;&�>���Eg-��x������z~��>�*�t�����0�"s�(V����^��8̮Q#>%���H3�ܿ�UརD[@4dD���ܓ��-�ft�o�u�
����V���e���w���렷L�,\ܔ��R��&W&uW�$��F&����R��)�׊�,��c�~�J#���X�Ǥ�ue T�x��d`a����I��%�m����d�[uSb�B=�3Y��L���,��Q��CQWY�T�1�0\����_�:��xS�쾯2($�x<���n��n���{-d$e�8%(h��d�aj�,�D9o��*D����l�v|��}�w�
kF��;���)Q��h��Z�fxM���_s�F�Մ�!#L��oA\��cJ~{�c�l���x+:E����Nov��ñ=V��t�)�X���r��
�V��ߞ���D��������H�;Ku�Ʈ�~��Mfc�c�@���N}ȣy���z��{�ӱ���3�2`��p�i���{�V��!��7p��y{�|�J_BBgU�m\��y>?����6"	���P��m|�f� 5w��A��E&U'L����^��H�j
���1;WK%�d_�R( ��kf2�[E�⫒¤莝��q['�ɔ��p��߻����?~9��P�-��,^�zo�� �b?}���h�%�+���\�v=�q��y |�A��3	M����7 ZҮ�ײ�I�5t�&e>�R ҵ(o/يq�5�bfR�l7�F�C�u��^®��X���ѧs��rB-�I��ƞܦF���텃&����2�ڊ}z�ޟ��'֕*f|�!��{�ۓ�ٔ��U���^���:���F��a/l.�{q~P����&N�}��q�?u�o��p���q)�h˽��
�_Ve5Q��ɗ�Rc�z��	�-3�f*�z]X�u�4^v�����#F�b��6���a��v�W{�7e�)*�j{�[[[��u'S��zHe���_�e�I�F��g� ��BX3(�m��iɡ�'���R��4N�;���1�]��3kJ�ۓ�Ҧ��T��n�g��q����H�ɉ���|s,�ܥ}a�%4�{��X����d�T���lo�rݶ��6��&�`P�k�#��8s�o��f��`�b-�)[�]��k��3Dc)SF'	�;���,���Z�0��$�{��LڝPXn�|��E���{/7DA4|N�vM�hUJ��,e�WV�K^�Xs���E���������u@�����Ppx��-���a����1
�w�i��Ħ����BZ�@�
:p|�k��>���w4���H�!���#��=#*l��� Jܙ^c��.AG��k����J0*,�\2 �G�`:@"5�b���ؑ�&$U��є�Ė���u+mg�Fj�1
�Oۨ_�����%MU?���$E�wd�`ֶ,�uR0
+Hϳ�%
��6~��e�|3T�x�Z�؄B;wK]���v����קJ1����P�f�� �Ml_�/�o�Uf^1��(bڃU/�o-�����j-�N��w�z�_vfz�*{?#%�N�vZ��S�Ķ������L�A'}Tt�6�=���_��N������YR�5|�N����0��nO@�(�}л%��MuN��ch{te�e��d�7�3��:I�h���0GU{�����kf�ؾEe����C�~�σM8](�������(q�)-�@:�{vm�9��q�]��x��1��c����L��X�U5�1�P�z܄v,����(�/t=�$���A��=����4�o>�]NA��a�x[�MR~�B\*Z�2���+��t$B�˵̎h��sz��n���
t�6e�:P���Z�[�t������z>v?�<�b2Z~A���`����樏
9h����^�����`���sg��½3B<>Q�p�>��|�E�aK�z��D~«�0?�$[�ZmQ�%��s����'tG-c�핳�j��%*�`�V�U#;��Nk1��Vjqƥ�N���,��~o�u"�Og�.�H�C����Y �s�Ҁ��1}ve2͕��aI�K�MׇM[/��̸&�Y����|��ߓ�s҉Qw�G����Q���柟dFX�
O+o6�ɿ7��(�j����;��촤��j9�� ��١7d�I�������$8�GKC���h�h�M;�F^�����c�Ё�8�֘�èx�vJ��>`���`���3���z��p��m%����G�U)-ԥ��� �pgqe�s�{K#���܌Ne����V���>���\�I��Iu�BF晟@}.�\f�q�L���F/e��v�����f'BV7�\���K3����X��y�p��]�Sf���D�\�m��!��
�Ei��:Ɨ!X�u���p�hҙ���2%��}�K��V�5K�`��C�����ݯ�
���[�T�b�� W�#3��n��!l�B]���@ h��i<I�EV`��X�u�y2v��p$'��}��n0܌�O�؄�f��|�+�Ea��1�b�Jz�d��_�ؕ�>o�z�p�k�*y-��!�=q�(�(��E��KSUen�6ۑ1�9�l�f�̔B>\m�0;�TmJ�?��Da��F�gGpנ�9��ſ-�L�I8M�H���%`�E�� �]G8;<^�V�9a&��j����Lah2��ٮݣ��w���Qgs�>��W��:x��ܾO{�[��ڥ���L@>�:�;���
A�=�xO�.}����?��d3x�!�0�zE�,نjr�V|b�#g��Q8������>��,,��`��E�(�h!L؃5ؠ>,���2U!��A,qi�|�F��""�H��Ѧ�"���'O(�t��w�W�0G����O��c`{JV���^-��Y#�}
�G���4��fw0�{y��CK��5h����=��E��(�',��^��-Λx��?̹-�]�IX��^m�oѳ�)
C	ћ/lGD��իa�vp��5!O6 '��u���uԵ�]��D�N� 9�H0^���3H:Ԡ�/�2^�M���b��K5?��$����MN��z�Is���e-�l��:?V~J�3�B�����o�W_e������9 ~��DWis.�Š]DH[/���h}@���r�3'�BBcJ4�Ҏ��̝�[J�����JJ�E�)���-��i1�CY׼;`�,�[S���OR�j�ߦd�\��tZ�)A�v��^�Y����%�����p�VM���wk�����X��Z�Ad������"��>�[!�������=��9+έRQw���#?�G*@HdǧHPU�h~��X-�G.()ʠN=��R�j��p:�T;��i	�کK���J���=�yZ��!���Ȳ�޾��ӖR�,��A��ԛ�R���)39���I- %��Z��QP;��v sx�d�@�.��ӊ|T��4cǊ7�������j��8�;����� $0����vΕ����:��y�֧G��4�i�r���T�J����?�|��|IԤ���Q�T{ߣ�k$D����O͒R�Ώ����Z���@t�]��ٷ�s�'�ئ�/M���N������н�^���"����^
2�13Q
����t�Єf�5����Z���`�<�xW	�({|���悎�1�ܪ+���*S��Z�J���D{�xK��i�SD��R��/e�}�郐���3�p���Ssk�:K{Hyq>�G��6d@�f��8����%���_����Aܗ���C��)�g����e� ����uyO�����a�E���7�)�^�8�reH[���7j��Ns�L��o��vn>��4��P�N~G�d�b�.�j��8fpH�X%q��X��h4ۈ��:""c�b.��x��c�5qx̎dI`}�	�,_�P��]W��d��`�p�����@�:QJ\H��� �z�`S.n=�si�4�X��
�xֱ�Ϯ�d�P���2�P܅�|��#;n�"�mi��;�o�2���2[��`/p狹�yOur��3
i���We�[�Xzf�	?���I�70�����dp�U���nj���t��k�'��q�ӈ�}�Sף�B�p� ���*4lǧRG,!�|���2����ں_�2Y�7R\7��'�Ie�gf�؄�y�47?b�Wmj���ؠؼ�t��)}Rp7�����.�P�Nd�Ċ4�� Zٰ�}\�
��x�"	~��i�N���Je��4���m��ö�e�h$�D��y$$���`�3i[�@���s]��'
X�y�D6����E Blx��V�����-$|�9Pz/c̸\��KV�0�!
�B�K��(��o�J��&`�rV�9�nf��s��׌�)MN�04z
|��OV�[`��٩uҘz�з�yTvH�!�08���5�(�$}j� �����!
P��Ψ�F�c�K���"�64��/��6���`�LS<kS9{��R<��z2��j���;�Ŕ�\�cT�.&�5�6�s-�:G���Af%i��`׀��蓊�J꒰4-��t���E�܋�8��X��G5�`/_��P�t�ja�V���"X��N��`C�Ѽ�{`�ϩN���|vy{Ci ���_7b�4�E���RU����ƮإjD6i��¾��vL��b�km���@~�����:F<���DÕ�Xn�@���|	d�%N��Ϣ �PM�	7^Db)ݚqHKj����~.!��S�7%�p��&�(f�=}���` ����:��� ��-���^U�ִωW�����3f*�z� �\�2��뵨p�戴E.���a{���t�(��wg�:��t��,�.p���.��I��9WAxÍ)��Y�����Ӎk�E���Z�Q-�{��:/�sb���ܙ����|2\�\+�*b�v�M~���{�`/�4��J�ra���@���9���%v��ѧ�]�H������=��G ���bʏ�9P�����Q_5ˉD5:"�N�O�?b_�hcNe1^��5_�õ�9n��#���n�-���i��OA�K��(6��Ub �jjHNΠ�c?��yȡH}3����n���b�U%�Y�0{P5s7O;y#"�[��ܐ_�-kS�˒�w�wE����HCE��=f����|��\�֢��d�e7-u��X�<t��W��[��>�b�^0��c��/$|�à��m����~9�Nl"Ӥ �FLx`�|n鋗��_�ԝ^OaFᵷG��Q��^�.�8���DW��"d����y�^��z��e��{i��P	�v�E]ٌ��r�d�j�0�o�<�0�n�A���A�<�q"�~��GB����z�T�i�����t]����YF^:���L5g4(�F�v�SE�2�}�q=F���*��N�w�LJGᗴs�I�T����%' �޼�)|2>�[h� I�>S�f��\A�l�7�m��!��u����'5�`��3eAgh���:쎹�`�'z��S�)���2��D����WF��χ7��4{ˇ]�;ڻ�����Yd|Z��-탔g&�VQ�������?���`=�| v{�m���(ԅN3A�q���r.�pə��2}}9��
ŷCl!�}D��s��H^q��Ǥ�*�9X�;��L�e���_U�]����Q*&;k�5�g	>����RhJ�����"���*�U4C��o2��99r#g�o�6O����*�TeR.-^R�>��t�/s]�#���yx�a��Ys�>����S��2�a8Ӟ4U��?�cp�u@l���1U`�D�#�kSX8:�9�l4Q��t!Q��ƶ�6���j��-^A���v��$�\�E?�:bU�={m�x��+{���|�,I�E=X���u�_3�����[G���sMM�4�O_Q���[L}��ȉ[����èO����q?^��<PKxy�J�j@Ԝ{l����%F�4֑^�N�ʌ����Yg
5��>�<�m�W(����ޛs��0H���=�I���� ^��q��+Ԣe�SN��ԅxϵ�$�3 $��Gw�Sq�!u�xk͉��y8r:!-���.�׼�
���n�r9b��1��BZ�v� '����}U��X�]��:C��v!�*i����IFʧ�CE�����D�q�K��TK03�u<��ó��:�=$4�DuH��.�Zaf�j1H.�S�^�W���,t#Z����} ��1��T���G�t�u��q=F�!]F�EN~}����	TpH��5��QU�z%9�o��#��56B�7�iD)��2k�Z/���|'�&��/�ka��V-\"��j�u��[�W�X�ZK������!~d�u�8�a\vlW�H6���FU�A�a��zqY�s����ë�K���x��8�e��:�<$��W�9�m柤��NQ�A���b�i�0��?Hܪ�EvѬ�V�� ����7|��	J�c��Jx�X��>pE#PJ*�Z7� ��G9;ˡ��4٣BQO��/�V`�k7,u3��p����J뀦�l����;ޏ<JT.�';�>b�q�<���k�ܺ�� ���0��N�2d	� $����a����5� v�����帯A�T�C�I��֘d$��<0(�H,���D�>h�[��=ϊ:m����8r���� �CC�*�7��pƞ��r��>6��.����-�E�a��	m	{�S���}���Zf)��&�t%52�$��-4��7ݬ^�[�H1�eg�郼�$$�#����&�*YP��?qO�M�?��VQ����3��=LAA�M�5ʍ��<���BB6?G捯�g����Q\�h4��	��Ȳ�%Oa�ve��ba�?D_Ko�P����3��ЪmcA]�Ո�k�`Ӑ�cuV�����W�}7���vҲ�P����fG5͛�>��:���á_(�+��KSl�H��i��Ǚ{�h5t�VSĻ�*���)��&A�pu�6�]����U0��VFW4q���(��ʸ�SR"�~�H�K���Ž���4Q_0� 7%eƄ+�@���`�Ј�{0).�),N��ԧ�U8E:5�cJh�%��NP6U�̣��Pyt���靧��w/8�-�����o���ߏ���\��%Hޘ%�?�-X�7�[���;���� sǷ�Y���h�͂e�����&Pz0nT��)����P�<�����_�*�]���^\D�l��9:T��	�'jm�#��䫙���w챢<���� ����I�A�k/�<��������c��P2D�^���մƩU}�w#�2 4������O��KI�Y�Z;9�:h ֞*�g�zw5Ri�9z�i����<�n�T���Z�&����}�d^�l�ݱа�c��1oWj�����Ev78�<8�	��H��z���EM�PR�-�c�䘨�os�����YK�����*�|B��t����]���o&� ��P6���{���r��Eξn�c��{���B���-�g�&/4��=�?w�\ �0DEX�O�W�ܣC�XМ�� �d����D�]�ܿߜQ�GS��&t��D���Kx3i,�j��p�y�Ĭ��_Y��E�!l\��)�t_�>�3��e�5�fB�
��0!��?G--�B��9(t��ҧ�q�:����M�܈[sXB��xKf�������>5Ě:��ڋ���\�!8�:��[����a./������j����`����{�����_�SV��@���׬� �|-�~3���Ne�ʯ	��s���|G��'���1�����.%�Fʢ�d��Sc����s.�#6��w`;�m���2KX3(�:f��=\�3��r ��=̛�B�֗�Y��K��i���2����60���"S�de@ʈu}�p���!��DT����%M_��9��bѽ�-X��5p�/��	���P�y��0݈��5�{�x٭��ua��6) Ge�W�{��3�b��r��+F�т�=����5���M"|�Bb-N'�X�g�{����6�h� �`E�D0��Y�`�c�Aъ�6���)7��m�F"�C���v׹�8�l��H��:sp>����/�MQ����φ���z?�7ɱ`��#��U������8�M�~�x^z��6JP'�o�CE��|���PJ s��<����\�֔6'�շ��V��=fCB.'��/z��1m!,5ĥ`�Lw�R
����n���W�-۞�d���a��ZvJ�ld��4�	-Gy�[�"(�ٜs��CA��'G.��#���xqOkZni9Ӟ[�1�=R��~dO�p�x�^"S�E0�,Ӊ��y�
z��x���v�Ir�c"8��va��(8�O�RdnH�IoOd�̩���jq-y %]544,��,/ub����{�0C+X���fCd�뉿�ir����Ɇ��F���&Z��]'s�=HeTx�/h�a~�A7�D�}�R���`�bWǢe<s���!��[(�*w�.��T�_�
��[MMꆳ#�d�����k,��O����}��R�ԙxI?�xW�.5M�4��¨�ʚ��BQ;I|��>�4��j��-�+y����׸0�g���	�+Vd�&}�`���ZH��,�=j�J X�0I���~�7y=
�\�#�MR��n�q>�PSg;ӂFenq*%!��FX�p���U+�%����ɞ�Mh�3��mZ�����-�7B�2~���!;�f
�F��Q�����7a� %4�)�_a����M!�1/�+��pJT&b󁫉[��s�x'�S�4�AҪ���E�~5�9!�v�ln�<� �/�c���E�t`�F����Q�mb�E؁z�r	��+զ�@�-P�y�&�*e�	U������<�̪7\��W�H��_n���woo҇���J<��Q�<p����k����'�y�Nܑ�q&X����ާ�j�#�jn�ҷv3�ɎjF�SQ���l�O���Q��'¤K�4W���[��P�N$p�!��P��cб�5�����3��\��f�����p�"�`�6|�r3���0����s�:���f)&	ߍ����ȋ!s�jҥ�~0A��'0���K��~;�Q�c���hRP8�_�(�!���go)�*�$�>b�.���w�);'�E�o�;��H1h(����|��1i#"��[�T3�To�K��8�	F�n��u�գ����� �kZ�+�+��'U�GAk,�%��̲p�z�&LSZ���H$�v?c�Q��P!��m=��hݕݩ�۽J��њ�r�v�E�� O��!�d�������9�a��iH���}���w2j���m 5i����+��ȗHyc�tP�}���'�d��^4\���_��Rz�X%#d��<�K�����6��ápk��E�޼h�#������8���i53�k����T���fO�����e1?l1��*T�e?�dOP*��0>�uA	Ë���0B�z��j���X
g�'��y�C��Gw&���ԯ������"I���TTΎ`]wm=�YEos������aK���b�$Z5{���`>E�u�ɕrv�t�(یf����p{�5&��&�#�mg������/C������t�̮�Dx��:}וֹ�DX;c��/o����I�d��S`�s7MJH�3fx�?UqL��J�K�Y����?4y�z�wkC| ��h����9�JN(fJ(ޅ-��D�$�[�n��w���2�|Zs�f�_�:���n�����8Vt��L�ȉ�	�n��k�d�C/"A��SY����f@��j���?aQ�J&��$2��D�A4�����-BB�	��6��R`�逆Ó1�vIy����'k�U���'�3���H���������s�G\*h�����m�������lO�^`t������1NX��h����N�gާN33����<hf����vЙ��\�y���ޅ���"B[H�b<[hG/�g}��s_�#�I{`<��i���g�V���\F6NG�����_��[�EV�ȶ�^P91.[l���=�%M}o�ԓ��ԕ� |����N�J<�{k�Z�F%�QDҋ��v������bs�Hd�,���ӄ���'IÛ�]N�=�*~��T��z����Ȓ�>w�D��k4�/��|��q�k� }M�t�NI�u@m�g����y��)0K�6���E��z��u�C|'�g�L9�F���eEW���uNq�[hl��f|�Q2��4T��o�J,��z�JC᫑�!ձ�H5\��D�6MUa'FG.�y���!}xc[G�,M
H����H�Cb	�@�;n�3��2��؀z�L�Ԓ1c<� ��Eu��y��2�zgN�V-W�I���r�/וWj�BU&��i�r��
�~�Wj���%|�����(υ)U����%E�Eش��*C|.�G�R�~c�㙑��n#;i��~��񏷵bC���K3�;���Y�4)UMQ�I��`Uuߚ`M��ݍ�S6q3���u��
Kc�YX���+�*��]<A]�P�e�C��:�?
%�fwH���8����n@�P�[R��<=���9b���|�k2W�aN�Pz�����S��h�M���BK/ �������i�2��7@�f����+u�0���I����W�|�|�l�+���;�Q��9��H��"��7���)��H��\]+��V)l*��k��쮞
�>�W6�	�)dF�SNc|���xG�X�����)��ٮ�X>v�^f&X������QuhnO�DIw&6�$B��a��"�r��(�c,�(��%�T,�\Ys��8חph2�C�aqD��3B����ջ<yJ�6�l�T��]�n+�1y�δ������i��Txh�;�#P\DZo75_�� k�#71(�ځ��#H�����'��l��>�yҖL����z��.�'�W��<+�@��kP�Q���X�e���I۵��dD��=���׳�Nl��=#��ƂF�Yx�IF����y�# �E���z.�>�Ms@e_����p0�E���t��B��:�Y�"Q�$��I�}ᶗ��C!�ʒ�9��[_��j6��Q2T��T8!
g���Ѿ9"�"��ky��g}�<H�p��b�����3�ne����Fl�U�z�D�����������s�x߼�@����}G�3�P�OMx�;�n��ѓn��� z��4����{�� ��W�X��,�AnV��BU���6��jS=���0�fxi<E����s����6��(s ��e�m"KE#F��[Χ4.������rp���j������q�������bO���ʨ�	w[����*䜃a�櫅�(�Ddo���IZ,�Yw�5j*�@3�e�(]��s���$6f�؜8��`5|oQ *�|�}\�vAS��M_s�o�~nZ?X�����S%w<�x���rN��d�2H|ϘsJ�ǁ(���u�1�^F�>��D�Y�|L"��rq��a����9ĜkX�d4e�S������@#��E|t���wV+ <H��s�\��uz8'���d��{X���"ʗ������B�h����{s��V�6�XV�sY>#�N�m�&�n��B���@>����솽��A[+ȍ��K�uy+��.�mH��m%��jN��?U��	��ܯgk�z����>y��Я˨tw��r�7�I)��L�u��03�,(K����鑑#�&���<	��GW���2�;Q�f��^`�$��!"���Y��jc��N,M�<�n�xD��,QO� =�g�����=���5Դۈ? ���4V[�*v���PUl�rD�[���0j��>h����0!�0?�2yB$3�"�h�J���U���ޟ�d�Pf�ㇼ���/]�8K���"�)?�fH�4�g�ם�6or�%,���Y�A��Ȁ�ę7���r�{���	�<�]Y����l)�O7r~�}ܲ�@��{�2?;������	���o�����m>�j�>�t�,f�~@U%M�DF�����C~n=�	�J�=A�8> 48ks�-�K��2��W�N���P�良5�~���^�<6f�����i�_i�-���rqz��0g�I/�Y��X����u����O��/`呂��^:��٨�홄�͙�=�d�T�V?��A��u��_g:� [1���x2�]~5Ƹ32�
C��$�E�)�t�3k[	Ծ�M��]�L�Ugl4��I:?��:���x!V��m2gK�c�!.S��H�(�ٍQ�1
�Q�!^�,ԣ�:���{��JY�;�$*�ˬ��ã�E��qw�/k03�GS�Z�z��v���B?a�u���az�I @��Y����Xbj~�몒,A�ȧtv�f��	+S��g N�_gNzN�,��v����N��^��<P�����8���&>p��|����u�V�3�II��P�J�M��}<����'2٣�|�n@�s�Oض��I��M��Ŕ����+w�GC��
������L���\���H�+����D:[�e�q%��'MF��L#�+P�a(�y�5�����w��K'J� (�[��g��U�܁ܱ�Hw`T�tU�rP���	��q$`������jh#�II�$ߛ|ګʏ�^=����!3��Al�e6�^M4�U@\�j:e�z����.�g$�o��/sd�}
�������]_{t}��
��fֻr����<N�Y�:�d�K�N�a�Y��җ��A&�.I�B6���D�����xf�y����	��]����F�6|�<B?��櫗������R��w�m��� 2A*C�+�q[Ճ0���0"#Cq���4�YV��=wH���l0h�h����-f�TP��Z)�?�篽O�~5-mF�y��3�����5C
& �q�&p��b���0��}�Đ_x��Y�0ڑ/M�,��*�:,� �����;n�!ߠx� �̖_���98蝇��5,�]�x/�ƶC��3w�4���yHB*H?m?���9�����=4v��[[/�jRMZ��>�HЌ���a&���,�}�$G_@ի���I@Y��ڱ�(��S�?@�~1�=⌔���U�#�ٲ�ko��kl���h�y� q��`�X���Ȅ�d��=uk��[����1���#/d�of}����+�j�#�S�$��~S��&�.��/03���C�p���^WM|�'��}.Jc�sh�2�� 쮁r8�j4��J��L���?�fm!����a�ɦ18t��Ͼi��6��	;�a�Y��~I������2��|��O<Ҽ��^��T�S����NvO�G�[�������N��4ZTF����2��T�-�_��"O΀)�j�=�(_���Һ$�^$N�F�ՋaSVX�.n|'@t/>^$3�>Ę�X�u0*�b���*�<���t��o�⯽�ެ�`��1�U�����Ax��_a�f���FYR��b�x��HD
6�}wO�?x0��6��r[r�^��.-���<tvW^ z�ϼ�)]E�Pwx���Z��ԍ�u����HH���g3���H��C6P?��$������u�C�,O����Z�N�]³��{9k�������P�د��ͷ�P�i���Nv�~�c����Vυ��4b�v%���[.�s�J:/���Ӥ�㦘�_�8.t�-��jz���x��H�4�o�aP�o�y����#c`D��0�@���s�hL�� ��o�-�V�Ju)��h�?NO_�
��\�{5W�>�IT�Kf�νٲi{��b����yj���.�!�e^el�<�ӷ�MǛ�r����.:��Q���B<��*=3~i���u��'Q6�+�v��������i�(�kۨ��q���McCj�N�"^p˦$�у��I`�.#�@�{�
\S�4n��~a#@�6^܄Ճ���#GR���c����z5#hGn*(����=��ު�&p�f�$��}B,�T�+u�mt�{�$Xp{m�d�:)d�?�x&Z�,H�eY�=6���ɐj�h)�F���}F�o�YϜ��ϱE���4&�]���?1\�5_'=�	4�A�_Vi��n�� �s�N�A���[�s�sa9g��	�C8LV)\t*�5Mѳ/ѥXg��ƕ7�ˏ�U5������P��%��=�")O�'�}6&(��a$��a����F���y�+��a��N�hI�\&���J��8S���Ec��A��m��y��\�C��b��=6X񀏊3��3�`FL+�qa'�����Cÿ7���^U�0��[��d�3�Z׵���7��K����E����Svp(0y���ͳ�T=+@),Jm ����`� ���fN'®�L�S��jY]��"��P��p6C[�' ��ҟ���9rۖ��Mk*ZaU��~'ty�I`;XG��f����=����c@hYg�`u͉���F���|�V�ǃ��r���m7�Wuv��X���F��
֪y@PmV���{���Z�(�;��7�g��Ajlz����M���SpEw Bb�vM��{M�8�_�z@�F���C{6�2�vf�F�ƮE����g�o �A��5�.EF}�U��p��S�Z�?��i*��;�"2��E�����i�>r"���(ŗ��A�ǹ.��W����Wlb�KBG�:���*b3�Љ��w�L��/D�]9e�br�OmJ���Ǽ=�쳨�غ�-���	����ry=ao_���!���g�!�ފ�U~�Qp���2<����!6[���V}j��: ���N�l�.%��|������,ѝƚ1r��db���JY���G����`-&�b�R娊ń�-�Z,�c[�z��!toMJ)i�Ļ�����'���8���c]�@��U`5/�;W��_�D����)_����;����yD�u#������@S]j�}����DQ�G<-����"^g��i,������#o����d���e[r=��~��{��۬�0����y�]-l�5�|S��>�LDh��7o���T���+��fiۜ�DD�$�/k�pD[�B8�U��1bQ\K�Hl~8U����?���NK����+9|�����*dr,'� #ؒ{P8;��-NxNȐ`��j��7��5F]-fǊ/O~{5}�����{�L���6,X1)�$J�5�iH?g�Lw`OӪQ�� >d/��tO���6�s���X]N.=՟äN�@e��q�����5�M������&'R3.������8�fS����Q�Y�-����i6M*�N�A�����#M\OT��i�=���R9�+�x�X��Z�N� i���4��G���1cQ��ѳ�E5ZF�ǚ~Q��I�A|��p�;�T�k�۹����D�:��b���jg�'��i)۾s٣���B!}
���H�濾���J\�c���"F5�k��Q��p���\�ʗ���	@lC嚗)ǝ��ES0�I>jQ�㬤���� ڥ;>zl�-a��8�L��u��2�dh2����$���6I@����aO��(_l0����c��R��i�����V�as�L�8`�Z�d��� &ńM����`	"�����Q�������t[~Y��&T`���N��qE+��y��Z��}p���x|�:����<�So����KAy�z�f'�Ӻߖk����lC
�6wڀɄ�1+ ��(�W���&��ض�;���/����`������N��Jr6P*���q;�R�>��3R#E���D=�����˿b�����+�sEE�U6�_f�㺿�q���*�"r�x��R��ZU��^3�m��P 4���C;Ӯc�P�^�U�e�6��Y��[C�x�+T<6X�q��}7$D�����y�ȕ���c�Koo�R̾��2����衱<���8_�@���*���50��z�+7�HhW\�7���6�oX�?�|�7m4��Z��컘5��ب<�w6Yg�p���r�L$��%������oD�h+2�ie�o��vb��q�n7<���N�n�Q�Ԑҡ�Sp�*���~i�(1�`� ��!�u0"�{�h����;NLL; r�����٪c��Ǘ�
�"���٘�9���B���`��� и�+��9Ō�q}�E/,��_8ꌝ�	�^5�^u4n1���VT�h��<�&2����R<N��*3��wv=5NR�����R�e�)�{g��N�t��h@O��#��QE�ݳ�701�J�sy�܄7@Մ��Le���M�s0o1R�$g:#��n$M��BL�$�G�]��ɨ ��+�1�a��i��֨�L��@f
[��Jc�
`��NB���cךc�3��R�H_v�054�uY����e����+��]�(�G��ӂ6�u��3@2�C^���YKPҷ{��9<w������)����-ohX���Sx|ZP�T/��&�&4�g �"����&*��6i��N�����)�~I!��Vx�dj���_%��NE�]�Hh�o���/(���(H~$����}2j9��Z�t@2�tS�P1��m�+q\חM~O?<W%�Qq��|[�k��U����a��I�z�$l��((���K�a5�c��<��s��N�#O�W��4��<���A��v�+ú��O:�����̣b�L��u ]�����qQ��<qG��J��թB r�i	.�eYjF��H_*�}o�Ȯk5�ܖö�0��`����.��͞� R��.̕Byڎ�^�I��;�Єz�W��P���6C��-5�ƃx8��Y�jΉ_~��?Ң�� ��Mr�r��ch��u$��h���G/=�#ď�'�T�PM�&\:�!�(_�f�e��Gw1���?���|R�ĭ^�6Ba\��98�C���$�@4<(#np���-<��*-�����|�qz��*��9L.e&�����3[9H�?���GN�L��� ��"6Qb�<-�x��f�|M��¥'���o�5sJ��́�%o����fR�4�5 �f���"�� C��Zm������ŊֆG��X�(�k��!�#UҀ��i}���*��ڒT�έ9�̓)bV*	�3fd��6�'��j-5�RI� �%`�j�04�5��W���$=��n/��o��Ֆ��Ez`���ɊɛB�\ڄ
�"��!Y���_���걪ܸ��9Դ�G�5kX��80�5T�r��(ۣ�������RjA���i ���[���^j��<�[���c's=�Qg�1�J*)�"��?��dG��L�+�!LZ�_���Ƞ	���ZOl�`G�0�d�˩[I���}Ԃj�Ϛ7Q���J��+��D{��)�%e�QE��J��!?*�WR|�ϯ�i�ÍUF��L�O�X?�Pށl:�L�>�w���ʳ~Ƣ~.��B�� ���LZ|]�CRB�.�O?�Bn��Y�c��Qb�u���6�2g^a��ܞ#�^T���
k<�����v�9n�A�ٓ��@�Cez~i�Dj4�,6�ގ&�g�Q�%S�hc)����lF�%�r`L�6[7Ss<����I�<�����>}�rM���\�#��W�]󆜧,���>Ҍ8S��O����nC�V3����}Ҿ-��h��Im���`�;�p�k	_���!1��Cũ��DxV�(k�zv[��c���st��թ�QP�z�MuI}��ZܥL5��`���.�[]J�?غ�x�~�v��'��U��1_��--�@�����z����:NW�%ۊ�>�K���6���T�}�3�X�G*��#�Z�������1�X�3��,�{��c�}��I^Y���x$���l�B����m&j��mĚ�H��5$Sb�B#o��d�b&�ɺ��oaY�ivG��-�@��ssf��P��S��%�\i�F�=G����{�1<�
2���@u�!~��p!r�xx�_@/�!{�9�m��.j�Mx���1��
�GI���:{ɿc8�5A=Wa�}�7J��6���4A�d�7�oZ��,�d��m,�?�O<�X/{�>��p4KĦ�l���g��k����6�o %5�3��|��ґ0L݆���>�� f�9���ձ=*��|�~�5���8!��04P��fX��UQ�q��<�Bd��_:٫ؓh��UE���X�q~�9�~},�iL�!�q��n���n�F�a�z?H��O�H�&g�����:���r�]���b��yb��у��!�W���O��*���1.���͎/�PX��N��]���4[���°�@A_/����H*�d�z7�7x��dE�p^�{�I��^��Z߻��:�V�ˌ�R�ŵV+\�ND��N�'@�]/`i7=�2#�7vȜa-S�f�����A)�j�d�=b�:�D��>���:lڌ$s�V���t� ��}ٸ����Iz�`�4���������Kx������(aClE!��\��9�����,(��)�Y":\�bo��n  �=j���g7����*T��a_案���Ҍ&k��MJ0���wx�oVMwl1e&��Ye�x��mLd p����֗
44%<�%��ח(<O]h������U{�"\��\��'�����Lk����7Is��=:�D������r�}�_P-l��=��n��گ��b��G4L��W�I�"oɖ: �v�[9WO�0y���ƻg	:nE�&/C_:���ǉ�h�C�b�}�Pa^4
�:^V�b�u��=�2���;'�~�������q��Orf�a+��)7wF�u&WG�A��v��@x[Z����m���K4���-]��,�5C�fG0����2r7*�bj��j���؇dO2`=�m7�m�>A\����p�ٸ�F�i\[�û�-G�8r�&SZL����N_��bV��tC �抝4xE�=Ri_o��Fp���e-�	�! ��׾����>2�p�?S���?eqIt�i-�4aO������������_�wWg�®~���2[BJoX�_I@�3,�#pF��>�.��)�1�e�۪��i.�H�-��zM��ɬ���G�W}�kBh���PR,����4�5p���E�+)9�q6V/�.9s�s��D�̵g./I# � ��*\g�xו�S.j�so��u��4[ܦ�#�4�/��.[<"� ���gi��{.�����L�1'	�?QR�?�z�m"ӂB��ڔkGT������K�L���--�D�O���P�z_7Ϊ�{�T�ڕ� �>���x���}2;Dr=�;b¬��K_0�!�-�h� _A�7��?���o�`EP��g�RU&|8U�$���W�N��o�D����xr�l�K@�}������_<���sKq����ze�m@�@00�LϦ=Bq�"��E͐�n=/	ֆz�Íen�
�{�� 0 zh|ß�.Em�B���A�e<I����J��lñY<s�A.(]�|&�q/�=/l��+m9"��h�X�.��>�VL�fc���TI�سR�ɅNctI:�YY($
�,�!�y'���1fX1��Z�m;���MĈ�-�νѓă�JSb2����f>ϥw6��>7խ^i��G.��l-E��u�lW��M<�����3��M5� Vw�)G�<3\xۉ�`��H�0�8���o~.7,�
m�]�y�ʗ���Qgp�����VH�2Ec /,�ǆAE����-5�LAcϝ��&����`󁕟��eF2��?���׆�˒�K0W�āQ�v!� %.�Q@im��J�ɀd���U���-�(��d�y�Wu.�Ž��>"#w�a�Vl[s=W@��gD������� s,��ỽ.s3�ϛ-�^�	�Dih��g����i>U~�
�EV�n�a���g�ᤌ8��ˆ����1�j9Ō�j�ȱ?������Ɂ��&�/�O4�����ьT�-�X,U���ܳWn>�A�7��Z��8~Qk��J�	�ޡ��u�ǥ��0PW<Ϥ��
w�����O���|�=�p�Xo�Ê3Ҥ��?�(
轼ƛ9����� ����V'��S4pv{E�M4h�wQ��k1A��:� 
����r2e���K^٠[��cj$�� J�e�:�M�kb���w*�>�TN/�Xh��/��]Q&��҈�Ԭx�f-����n�Hf�'�e���-.I&�K�Z�@#7�z������ �"o,0z#`�D`{�N��>˂�p�Y0?����6���d�A�qՕ껺�K�
���8ٌI�_����W�aA��]\�/������;�^A��+JR�RՒ"Z	���D��za�ێAMv���u���x�E�5��J��.l�@�8�r�����V�$�#��4t��zq�F�8��?��)ڷN.J�6���Nrܚ޸�M!Hh�f.���%M�*.�Ke>�RRmO���Bx{��v]u�Ѿ�+K=�FwVЪˎ6h�;��OE�������(i:]	ӂo��H���1Ƥ́��[� �NzȖ\�)RZ,m!�{Mhz�^�J��;����+�6]�ԡsE�x�E�x�e�����z�
���;  ���X��Z֙ho/_n�{���@uG�Bpv��(xF��*�"������uD��q-�o�i|�i+�WEMh� a�G�.�֡^�&W�z�(8-m��b&B��K%,�n��z�A�5'N���ӝs�!� }J}:GN6�{�߹T��;I���y��R�)����\eݵ;w�4mY����G�-��؏�_�5=�������8���2��S��R)�W� D�$7:XK�}#s-�˵��X�+�U�B.�c0�%1��=�&ql&�O<ߦ�U��ѴKE虫���=����]'����jƁ׈/�u��Κ�~�����ȅR��GH�G��:�	�/밦�48Ӏhw���Z��:��dkD�(�����K��hޏ����~�l�#gcD����;4�y8�>��"�t-�3�t[���o U
z�� (<lr��AG=].F���F�7_Jl�q;Imqѽ��ϪcT�L5R����/������r��"��G�L�s4Sg^��e��Qt�sK����A�j�,X�6IE�$Lx9���4�g1t/�L��6�3z�����[����e4Z%j�(4��6;�����b܏�W��ZIa�5q��x�������?���@P��3܂R,�ܢ�%9�/_5 &����?�k^� ��C5�9+v}�}�Sr�5�=��Pa�Ր�L��lcΏ��(2���%K�`�p��S��4�m��j1\���>�o��u�ԉ]]o1L���tέ��WM�yBu�y��kи]���ƭ(�A�W��-�z�b�s/�r��j'8�OңzN�D�:�^+A����u�5 #:�7�.pbFK��쁄���� ޲�?���"�(�*�{�^��̣Hv��K6���݇��z�m<������+�+�鏽�n~������n���g�$�}�i�mڌ='�X�����f�Ŏ!֢m�N!�9��J�l������*��uP�w�\�򎕠e��(��rjV���P
�@�ިu�Q���&_ev(7���P�:"�T���n�82uaA蘧��$1��J�J'YA�%�
�ɂ˪3�TS޸E�Hۍ��ټY����ȣ����VU��+��o��f&��������oT���-�+�[l�s�_t��v��{m]4.kǙX���v4���/�%u�+�y-y��k��Z��e�,��2�)��������,Ò��JRL⧰��@d��R�u�R��enù���l��_��P~?.6x�~�'��9D�����m���.���`�ck�I��&����e��׾V���@�|���B�ǩ[��G.�� �O�{D����a��1b��}�m�����x����*�w�Ҥ�o|Qj���q�?���X��eP�߳]�[�������:��N���k:ڿ�g�1Ȼ�^����[jƾ J#�%��>��yu�ه�p�L�_��?�)����w���n�'q�%�Z���_I�AM������rdT �4	�f�W��h1����|�I�wf@��%�d����n�em�%'ߪ9�Y�"PS�MN��,��υ��y7�Ą�[��g���Ԛ:&T{{��5q
q�6�V�x6�y�d%
�f�'�:>v���DsG���ƫ������ﰸ|��K�S��l�d��+1j���*�A�Z҆���$m-���T�bR�g������/�E��3��wD}\��Ҥ�j�S�[�}�`���U�v�)���V�2,^5�W�KS
��M졗FB��W̶e`t1u�˖�h�kS��- ���mxe��#�<4Q��������v��g(	�c�O���c�0Ho�m; �D3AI�)�� ���UT�͉m�^��Nz�"�=�t$nd"L�^g��� �Y�E86�{�.79,޼�H3[�������3�~	27	���Eq~[�X�\�qn�	���0g��+W�ִ��������Hk����Yԣ��B�I����>͜����~aV7�ÃgR���	:��҈=�8�]I��3�T���v�`��ڌ�3fdp0Nn��d�f8�`����Q�ȁ$p��X��}حËaK��iz�_Q?��(4�ɰ1�܂��0���V�)���+ß]��<Ty���V�*X�a��B�^d�D��w7!��T��*���m�D��kUo��\O���¸��Ti�J߶�wzF��~̀NN0�:t��TZ��X7](_���Rc�e���-SyPi_C'}|Ub���T�7�e�fbD�cG;����Yzhv�����6�5���ٞ�R���f5����l\�����4#����v�~g� �U����\� �|}S|������?oZ�W����J�ܜ���7�a�b������)�B�X;���ǹJ��qVN4o�&ic�k��fe<@~w�T��M�QB&�>_��@�'В�?}�.'?J��(�>l���T��4;�z��������-@ÌF2�a�1���_W���OB,a	re�������U�#e��l�#/�����	>�g}��LQb@��E7���a-���ij��[+Q�����
��䤫����wi�L��������(Gd.�^3�6��RWO����py��A��ۊb�R���E��*[=j��hP`������XD�Ju�����A
�ϸ�s
'MG�[�z%��ݬ{����gto�V�:o{Mm��tJ������Qf�o�A�T�cN�q����ig�Jt�b;�cV-ArX��mC6�&x`8#`f�S�����U�O�*�1m`�+y�z�F��O>3�z����BVڹ����˿k50�F�!��\�qs���]nK.�Y_-�q�xC͓��d��ͮﱈ&H����Q�?	�-����	����^B劗ݚ~�!X�@�zBC-s	Й́��t��u�L^�.*�{��z�켗��͂�0��֛��/_WG��Ǿ�W�l��h���?HD0�
��A��-�=,�Ql���K2#�',�Gx�^���֦FU<)�?h{W�An�pl�b$c�F����B��G<��:�u�n�'����f}��&-�@��{c{Q3�,�يE���0����*֥��?YoT���^s�����ͼ9ۑa�Wa��e�Hm0��|�s�>���e�s�J#���jʃ(��q������υ0%�=�fy@�X��"I��mX��
M8���#9t�$���_ȉ��z���
�ꚤw�j�����8Y��2�rs����"Am���##��)��g���5pڬ'�V&.J<(5��]�����%�¾���:F�s�l��)��ٍ�o�`�HU�b7����%��+ԕ�ly�"K���o��-���dR���=ZP椛����㹬�?�x)�q>�4���B��6���<P��p��� Ki��%�Av����*�D֌�oVc�v���^��� tC��if�%�2�(^dY�L�55oG�m��4��;.�m���^�i�6,O
�ca�͆�چO���>��c��=�(���	
�5�/ݣE�/�Jc/J���A<zᰭ�����ߔH�c6Q��L�oEC��Z}�f$|��!��8̓�@���Ɉ�A�po��z����x����T�	��!�_,RU8��`����W�ְ`휢�K�����:�^�)���� 	P�5�,[OuH��{��ޖ?n��E��Y�YS�'��R匼nؒ��fE�n>3�o��!o9��ք����f����uL�B&�נ��+7}3^d4��W�"�-Ϛ�M�d���E�X���M
�|'��/?!�t����"p�F��k�O�C�+����6�t�Ԟ&�"�{ɻ�7t�*�t��=r����`۫��z��B�������iR�����+�/'��_�l6�����V�CSږʋ��[��Ѿ���du�*E?B��������tٱˀ|} ���o���M��H�HX���A�%���3W)�~	�J���4�Z���;cB�o�*�Wl���g薭1�Om�>�>���p����#Z<NP��p��U��	�����>�b7^�GaA��q��`�k7����:����X�֙�?
v{j�'������I���/;��(������
h B� � �-�^o*���������p�*L�3�1�ȩ��1R� ��Q��6F,֨��ݞj+�S�6�#����f�hQII'�R71��_�t�����4:- dȮ�8�H��H���e55��_��`�Z�ܘ�i=	PTm:�qY8@^�ɒN��9�n!��6�16Q>r�ˎ�ԕq+f�i�nU�F�������d�+�����%�Ҭ��H��.(��eG�]�go�D��j��W�A��m-o�3*��9_�Ў��u�b�][POO����(�A��kr������R0�D�����Fn�o�^B°��0Ҟ]P~fǫ��X��$\��c�T�޽qn>��y�,M;�/i-���Frr��UcU�&�7O8��f]sK7b/yT`�A�u	�KT�Hb���ӻP%�s|C
񼼄9�U_�X�a]���ab7��E/C׉!hT��9�������
OiB�*����X�F�'�\�)J8D?S�Ќܠ۶N��bqķ��\ڥ����Q�N'�W��������RX)�kV[E_��A�ݯk��O��3�{�� ���6'=�'B�(�?"	JB��W�����>��1Jd� 	�Q+=���G��a���V/�w^֯mq��7 _��P�z�SH���@&��U�U�-ק���_�����ob{d�_x��NPu���f#b+�2��\]�uw@~�xD��g�0v��NӠ�s�`���ջ
|����l���[
�Wy%@��F Yԛ������ڍ$���:e_���1Ƶ�;���� `���N�?}�ms���>�T1#R�� B�] �&9�0��7�p ����j��5Y �j��
�qq��|ݐ��d�FU�9�'�'m�~	;U.�n"�{�P
��@$��4!5L����L�Pe �[�<��F�?1��fﱎ��[�*��(���f�ߙ�"�A�OmG�#��!4��ދ��C�L������E�/��5�����&��y�:}��E�kc����s���K�T���Q,���2L���ǒ��9A-7�v/��#r�#�A,aФ�}�/�q��k\�����i��9��7䙍�d�Q�ң~�QźJȢ�)x5P�;����V�68�`7�*R��Y����d%��o���Ɯ��lV#ӻ�g��#��A������In�ť�1����+�ϟZ?��I�����:�-���M?�z4t�x�@@��׀�]�]Y7���x�*Φ�3���������m	��p���?5�������#׹j�r#׫��Nz��� u� �9�/��n��MR\����d&	�8ܜ*���._׷��6π3X1�N�ͯ,�\�ˍ*�ħ�Ố��7?3!-9	��qЕE�\�9�Д����)�|YRtH��x�fF1-���R��eK�%��D*��e;����Jc�q^��B��9���B�X��M�:a��@^iP��qd�P����$�d�_|��N��YB>�~ٙK-|Gf�k��q]+.�~}FR��U�>.!ޝ�
��$>�QA�A|����J�Q7/�oG��S�3��S�[�©�JA��*
���|N�0�޸p޲1*u���5vD��|Pw&������YM�F<|��?E���V�_��ju;�'e�|y�C��Z?�Mo�Z���rb�۠H�o���"t�|�c|cOgy�7�k**�렩a(�i�?��:�!�É�4�8��[xW�O�]�g�n��e�+�MԸ������1��>�0 U����d'�!�P�����$�	*�oʴm��:A&��x4��X���O�1�Mh���)�B��PPR���>�}���Eс��,
����!�L0j�L΂f^0����T ΑW&V�4��������2���ϻ5���8(y&(�U��|&�����߉aQ���B���z0'kÞ�8f���m����䙥����\%ʩ�/�	Z�Z�gm�yT���ߛ�|���p�t��c�-%hg(�j�昇\J#cR�D��� ��@�s�w$�����3����;��3�DˑĐ�X,��U���d�$3\w #�3b�>��b%�4>po�s�M�j���*cE"�CWc~?�Ԛk6.0�N�H��T��?����XO�T(�U�4����B��L3��V��h@�3/F�_�v�:c��>lvcOt
QR:2� ���Λ�i/�Bf��#E߻�N�n��h�K����@��pj�1=�JA��!�P��/����������8���OkLx��Xp�3�ޢ�p�A���n��E�/y#��f�����2q4xs	<}A���@�������>Z�y���=7����Y]�I�1T���"�%{&1�҇r�3�����@�t?��q_���XC@rU6���Y0�j�{@7bf4�zJǪvJ��?����n����f:��St��kF�7E��Ń���N�/���c	8<�㑔�V2�u��M�9�}�����_i�ّ�����x`?��.�C'�hk0㍾����&�rL�Cc�ǨrR��O=�����8�'$.���W�p.�h�������u�"}jb������o��\Wp������c��V�e`��+�E��h�
-ӧ~�Y+}w-f��M��j�WǪ�c�e�1	,����5�A��2���_|�k���8�����춴H�okK�t�hi�m�av���9���.��7#�&Υ�]�S��g��O����w�7p�ci�sս��(���{ #*�9�1���������*~�l�� �S+���\�:B��`k�KL4�{}���̥a
�z���V�Po�.զ�{aX�Ob㚯;;�q�ԧ�g+��H>*e�o��H���c�C�^���V�D��J��1��b�LA$,�`ǰ݁��R�QØ�ZQK�<��Ѓ�*L�j�A ��������N�nagF�:���깛MH�@��T��K�X,�ߥ���W��������#�ɭX�%��TV���3�\洜Dls������e�TE��h3o�u_�y@5�J�i�p!��k;���x1P���3yD�c=��|7��+�٠
�?�� r$��������+ooװ
ŵΥ�&�U��N,�@XI��#4}���MEu$�^�&�,��1�H�j��6k�.���K�W����o�>&��]��$�}�$_!sJZc��ʛv�M����cbH��[ؙE��/9�����a�_���xg^�*����N��~�������bh7dB
՗͆�LT�'�w�����q{\��+݊��(Xn�uիSQ?�S�U��"kd>�/u�B���]�sE�V���Tƽ˺zG~eBrS�; ���y7�٧�s��IPK� ��*_�{@�}lP\����ZvoG�𔒼g��vL�esR�k��z񰯋��ٰEi���*ㇲ9�	��������-g��6B?�������jm���z&ߐ�'DQ,�� ��6�C�ȇ�?���v"0���%~�p (V�![�X6��9�Ȟ�&d��v�[�E�����bt����4��#:�'��d݃w���� c�v���uQ��dpx�����4���jo/Q�%��p�3 ��G	=����ܖ?TOL��0���,�^�[˱c�Rc��[c��Πo�X��0�ʷI����a�:���kS�w+�B��4	���#��v7�iW%���ꁃ����(o]�SW�R���4U��[�4��փPN�=i�;<}�Hٷ�ݼ��7�l��pɾ3VY��Lc�fI����� �Τh��-V��5�.���y%Rk����:Jȱ���`�h!�4h�9ll����2M�������e4p�7�*S:��貃y݀�a�>N���]s���ۂ�'!��!������Wm |a���^g�� ���t.�V��Ī��KS�����a:%
����bx�[�2���H�OHjC����z��gr��7LF�G�$��/��>�0f���/C�kS��')���!V~3�������|��+3��[�|t��Ao?��4A�D���gQ���⌀=��ċK�u��Ex)�	��V��!�.�������K���L��=��5�6z<�C��}У�u��2c����W�Ĳ؋��kM�3�Q�C�9@�-l��*�F��܃�(1�3�V<�4��h5���}�#�T񔐃\�\^�WR�B����#L�q;���~;��ֻ��uU�}�f��4�S}�����ٽ8Ē�T����,L�I��WЦ�C����G'x�dF�?��~6g��6�3G_�U���@)�����-�R�(�!�U3s�}[�Wvr�j��y�uT��S����+��È��R�Cr���7֘���`Q�� �d����\�4E6[YN��٘K�hB�0R�N���c������ �l����0z/%����RLt�	�
��e�Ԝ�<��vQ�.��,�I��߈�{���Ƃ���oB��5��ex)���ӭ/�`�<�U���� �&/%&�<>m�
��h2=3���+B-��א�][fZ�yh��u�4�"G��H���ܣ� �B4|hFo�S>�$*��H�f ]j5�-��;��p�R@��8�0�d�>��c������ �K�y,ю�C�&����������*���)>AY�v?�d�)ɩ�:�L���~�qJ&�@��Q���ob������n|�(T��pСW�N�z�	��Bx�u0"d�3q>�]������H^#�c\�*�jT�ߛh:�w��ٺ<W�ĐV�����D��5+�k�}�;�nL"�~��u��(�r^
�������~vt�{���6��Y7g�.���3w�	�}9�ᆆ�d3Dr1�����\��hJ"������+���)�M�g���T�m�`#	i��PIi6 l�^�9XH�e�-��Zf��fbS�;��j�5�d�N�;�L��]�\���?�-E�Ղ崯�
_��L�xg[E��f������: ��u�e�I���
%�����#�p@Ž!{��5�)��lI�竫�����CT��X�4����3��p��������OR��u�Q-I@M���?)$�&�?\�2Vw�'a�Z0;��k�*Ba�J�uݲ(���U���2�j1Q+t!1�l�9X���u�Y`������3}h-?=(iG&_�a������B�
��̌g�=����*�Y�#�:/��"fs�B��Щ��:�X��
p:�uw�ZΥy�A�~��ܳT,��������kT���t,��ǜ�j�5;�S���34!C�,Iu+L�!�K�E�&S.�8L�XL9�(�,��$���X9��eͩJtO����a�'"/i͍[ب���1��i|.嬏�m�jce趰�����,��w���R����A٦0�t����-4C1��0ֈʙ�|-?��sqj��m밤_Z�G91���JP����V�O&f�_7ֈ �p"A�@}�yXf��?	�Lg����Q�M�}�OH�툗��7�c��h`JD^k*����nЌp���O��Fٛ�b,�яW�k^�G�^y/�[H��NbLEht-�*"�	��/��Y&V�_@���Eh�T���������6�y IV�xKX8/.��q��i�����P�ʵ�Y��K�~���[��[����G�?J�A�����Eκ�h[\���(oܦ��,P;�vA o����ؤP�!��^Oڙ�� �?,4�&�V�D��3��]��v�|�:P�5V��A#=�j�v����:�i�˷5��븲vl��{��󴐱���]/�Ti��R`��<�q&pPbmO���ՠ�ѱ�ȏ �N}K�ύ�q����ϱi�9�af�v9�S���(d���.Km�I4�1Iκ\ɓ�-��-��&��&���lo��	�����ѷ����m��B�qcI7hx��ǟP\�]-��Q W^R�]�2�O��2�#WJ�!`pI���<ܝ��z�����W��uF`nl@�G)�+�&)��ۅX27Z�X��>�Rj�;��kQ��z�x��`�.��+��<�`�<x�Ա���N��[Ny�Q�A�Q���H�����T#%�]M�q-r�>��^�n�ش��O$�)% w_a
;w�^�N�`b�zĥi���w�S�����u�~<&{i��&\t����G��L��ا
|���v���lZ{T&ڄ@ˢz�o  7�p>g��퓍���9���b�Cd'@�l1��k|¤���^PiF�~���HG��� i������گ�bu:)2l,2~�O�vg;� �Uo��~½͓����Ez<*���'�
v��t���&c�K�Ld��# _�S{�r;�z�t��Ơio���堨홌�@�@]>���	��Q�8?�������zT%��d��ܣj�Id5|a�{$5n6� /��R.�#����-ي��D��G2���J��6�^h�ka���V\�ʽ�pW��ղKC��}B
���(.�RLa
5�\� <�z�rp3߮ �����x+���lh���9�Y' ����>��M@BGdŧ5 ���%t%�'�g�s�(�W�����;��{���G2 OĄ��z�JK����Jlr?Zɏ�����K�V)��N�GiJ�����A���M�M��V�Y��x��ڴ`O �����1RJ�淅��7*�#w�89�g�~����m��0:G=D^,'9U��o�������v���F�����SM��v��7u'����YH��~�0�z�#���ƪEӠ����(���T�5\�g*�I:����罿�k��J�*�B���CF�Pft�Fp����_!���y������f�,��]z@�3�����$w�Z߫�9�H;�l<w���X��#�0~���oh�B�j'k��8��2��@^l3�2�k<�����K��2�9 �c���qc�U��X�@f����=�b���@0��R@%
�"�kN�	sf�OEy�>A`��	����8��
aJx��	E���1J�re��V�� ��y�����!�!�C��	J{���\���3���G����BL���sBu�sV��^Q�o����������[x�WL3�I�PEҐ_���	��#( R��{���l4y{k!87��@*�����nQ�4�Yh/ōg�j�M�z���h�Pb`��Xp3�*TO�vN��ގ�k= �'"'���.�]��1�lg3ch�VA�dy�Q���eW��'AV��p�J�? �*�^|��8M��(i7�R�G�����A� ��e��8�}���^����?�ps]�O
a��֙CW^�'�#T���gC<=x9�Q8Z1�s����J��SZws�^C��q��D>Md	mF�%WI��&ev�����]U������܃�d�PB�w���6���&�#m뇛NXcmg�b�0?P���!�3=�Y�X��|,�� ǧ�WyB�m�ƞ�5��-o]CNҺ��[��ڠ��	����->�f]�Aˆ4��;���`�Օ��읶���1�qA�b��!ɠ�==�*Y�Ҥ���2:]]������}��]�W*��dy^�A�H�6�R%,�	b�S�~����ǈ��jy�,�G&.��B	E!�6�e>�MDn-N,�+�[A�x�V0��m7�H���b�PL�� 0:PzxZ���:+S���J���$�d���n�7O���-�q6�|ؠ�y��5!�.T�Ҥ��)������J9�4J�GK��0��5r=ܔ�ODQ���|��ѡ�*S�U���­&�.�O� N��Br^M�C���k�'�SB���
��dw�"�*�j�#s�����>Hcƫ��^�uCk/z�uP$D�W�wyhJ��'XQ%�ڪ{:s��2U<!3�(���N�Zhy�k&Cep�۠9x.*�(���1�5����ι:����Pb]I�ʖ/�6O	�y�/��Ɇ�?p���mҶ��9N�.��~Z �#i$_�2u^�Y�7ĩ$wf�#y�z�+�Z;�q+�d&Nb�J=���]�+�'�i�1��Ұ9X[c4�F������*,�#�V��m툿wAo�h�a��3U��ș�Ed9��|����l�Gl���8�5mU帡xq����A�*J\〵|�T�Cv�=",�X�T�N$=.L"p���k�*z�t�k��p������S����J{�|�����嚿#�0�E�!�	�J�t.����/�[q�� ��zh4#����q�g�Ev�%0jJ�!���Y����\�<閘qƽ$,�29�I�Y�$�����v�~o(�Q����#������w0��+��1>v��y��a��84Л���w��K�L���ʎ�������K@8��Y��sv;K��s�{z3m�1�l'Š��D lF�v,j�rf���S�*��(X�f꾧�oa� ���
y�\Ijcԉ�ɞ����߰�1�]1�$s�Uѭ
&����U��F��s�ɐ49DGJ<�$�W�3ܝF��XuP����}1{�2��R�&���#�7��
s̈́�6��cog���4u2�v2.�Kx��'��.���x���U���K��;
G�_6�!R�c~�Ôzbrb��S�e�G�����B���W����i`�˴|���	xW����;��o�A��|8ٙXO�W#�<�VP����de#�ʛD��`��k�� ���Z�{t�ޘ�H���T�����\a}��꿸�Eˎ�5�5�m��ܴ8����9�$S�vq��'GoKc�Ëc��h]�D�ɨ��?2�����=���~�k�\6�k��J.�Ɨ7=��c�K�n��g�,����b�$��ݻCO�.x����J�e�f"}�����ӉO��$I�O}�� ՂS0��
�R!B�Y��3����W)#rYS7�bI���d�M��[�Co��<g��C��%����m#��o���v�İ���E�(F�k�>'1�a�T��88!n9�N=�B7����[qㆋ�������F�}�˩�%O2�Cd��rJ�p]�p]�
���������Mr2R=$
��Ȓ�-nF^��[�h<���0pH�ϓ�k��QI�O��L=������T��Dٔ�C�`��S���	W��:���-Z��?w�l�}���5��5F�A]r�5�.e����T����|έO��n���?���g��p��u���m�0���*DrE�и���2՜o��qׇ�L��3=ƀ���C�5{�E��.�|R���j��)���r��c��)k�����4� ��h}W�>��^7JY��h9�鱙I�g�~��Q����������S] �����CK_/��Zz
�Ă���Ju@F `nt������h�J_bE99�X��	S��G��o�/m^{�	�:����CKcf����ȋ��T�8��9>M��4$��d�5�!�
�|��	��6/��|W�����kH��B�G]��i:��W?�7U���M��b��'������;���2y4�V��A���ƿ�8D1'�V��.\�+g_v�S ����k���K9G��#���Z���H��
'�OYb�a�I^��J�,j��G�o��ǀoy0U�R�*���U �����pьѨ�@�"���Yt��[� ������~��F\�	�4{�]�M�5kô�|w*Zy���O�}�_-�*5��[!����Ջ]\�Y��{��m�fe'Kf阃1��8vj�'�\�>���/��:��%WOQS;L���Д��u��v���h���9^<-t��$j�PxJu
�YG�BϠ���uY�*G=�ݕW��E$Ƈx�ru�Hl>X=�4/�i�o6���5�]nO~#F��j����u|��GR�\�mOCrɵDR�>o1S��1���Kv\v�J�)��4�&A>�FW5&j�4�1�ذ��1*N�7������/gQP�p�����`&4�cnJ��7?礙��o�M(�mR5�-��6�XۓH^�����UG��D��D0W+Q�dL������ �`�h�K
!�qYџ�ٳ�h�G�,�����_�w�MG�a���r >��h"��2�W��������n�R:���f�K����xd��Cͷ]�[<3n��x�ђi���o��1��h\�����=�Ͷ���W<�e��pk�P�]��-��[�F�'����)_�g���_��]gr�"���G��5�����3�l���9��u�ri��Z}�(�x�z�-{E��hO@�tR��D��;Z澛??S��r=#�jgl��ͥ�$��H�[�_�V��#-}X�)����f�F\rr�?���>��+�?f���D�nX�h����<,&�I诠�kH���N��y�6��Fm��]o��� ��}��-B�D����};�O���#�X�P?������)������h.����(=��v� i9�)e�3���ߤ���8CKu�|x�5�K�x�B�����F���.<4�m ��;]%����ӎ4|�k%NY^r@q���x�I㕼,lIA�g�����w��wt��i�t��J�"g��,?��y%�o0�g3v�
��.�#�Q�ݯAz1��dm���沅����31�C������^�Gx\�h�쇣��N�Eu��٩�䃕���EɌ����O��w!���9�����T��Μ�(#{���<���ז��G��hG@o h��
'H�ә���\9^��$�z6��	g}v.���nr�v�q��f�X7��^F��k��i!f�����ys��4.��P��u~�H]?צm/0:��+��	YJ	�����a��e6�����ݔ��pgj���@{q�-��Z��)���<߳p%7�֔3d����e��n>�~ˍ��u�kkW��?W���˽Ď�M;[S�r��R�����n������W~��z�R��b�Q�p�/��W�=�����V�"@��cP�|c�R�N%vG�3���]�-�!���G�oJ,;��U0M:�i�ޯ���1�8�8ޯ�}S�C�-�j)7��u+�K{o��c葩���ly�Mv�eg��
�*���-��@'�Q�t�#.s$؏�I�E�O~���'k/Hܔ!�j�T���BQ�F�(=��@.���bj�W�px;9�idW���*E��Ů�x���t���S����4mD/�}�5��>lG��N^��@B���,�C�W��dU~ZԚ���Bq���&t����Z�l��O������Fg!7p;��/����Oȣ ���៻��%/���I!V�!ႥF��������%- ��v�5�JC���v��T����&�FZ/,�ﻐ]=�x�=qO2@.��Oj�I����,y}�Vz�-i�$�XD�-Vm�N[p��b_Q���Ƣ����s�����Ü@AM�x�Oo\C�����i|k�g�oջf�����V�>gbKķ=�Y��1;$R��d0+e��/���\%�Y4=��aT��9�i(�I�Q_(k]q��pPh��T燾�̪���H�����s���L���16�F_G��B�B��k5|<w�����̸ ��X	RP�h���7a�a��U�4�}M��{�.��)C�5�@x���G�	&�8tI�����R/�!�c3�Y�T��R�J��B��_�c�q��=r4I��*��h�\�1\��t���s�a�6���W�>_���DR���\R<��-��G�1�nV���Š���fs�3�U	���iP�g͘;�[�.���s��)��D@�����bu�,�T�v6�m׮"�wp�S�`���G�a��Jb(�
5���6��&�h�`>x��2@����i�Q�U�kƉ~�w����ZzԓӖ�K�j33Lk�b��fXS;w%����UXu����v�6q1e��j�h�%O]����ƊF�+ɋ*E�=ق��(�;-U�8����|�}��3�\��MUL���,��G��N,5v$=3o����;�Y�ɻd��r�V���U�?;�s��1�z6��TӇ�"�~�q'�)��yS+��amZ^^ K8����n�gl�c�tz������}ď#��}7�o?4�T\Xw�b�~�#�w��&����	�x�O��g�3�ow������&�S������;�cn��P�����<?�X	Ռ�8N�����QF!d��	��j���X�AD>ů9�J��L颦�c	�뻬�[b�l����'�x������ft�N��ۈq�%L�Q��F�v泲߀�\��Y:�4�"X
������$~'�.J���bT�2C�]��g��ZL˕�S�|,b=N���&qMy�� 3_|3�K�w O����w��Q�t��.>)L�����8I�͈��9����a���!��StM.�挀�\)�D+'z��۶cMW��%,|�R��FI��}+5�x���p�'��U�0逾�ɕz���3���Gbԏ�}�<�z6t�:>�
�Dr��*?7R�u	��9I�f��υ�F�vȜD�үZ��)XQy2����U�$�����c�րoh<��N�����#����Ae�'#���aQ�P7!io'�z���Hw�;)E�.�:�-�,���|���_|��N�Ē�|�fG �߼�ik�B�e�|��?k��%��/i�"g^a���Up�m4��*�|j���� �C�<ҿԽH�ђ�1�����K1�sH�`�K�����/�t�i��`��1άo?�NB9����M̱x�]�$�/��^�h~'�%��.!zЖ4ߜ��ri:�8s橨� �8���_i���=:j�����W�ZO��w�ƉF�6�rhl��0"��iSa]�7�P��K�A6v��Ĵ{�b�o�j�nr�kV��L����f�1�J!4V����e�}:<o(C�S�����kj/ըx}Q\dI���s��
CEʚ3��vM�M����;���XЦUKDG]�R�%������02��.�=��N+?�f�0 k�ݲ��:��Xǒ5���1^N�����LcG�"	q�|>f�Κ�ц��{G���\��fJB!�km_����e�,���cY�eT��YxE,�����J4w<�s�~Q�ϾoK��v������n�a�Mx?�����$�/�n �~7���|�  X{3l�Tsie������Yd/�'����=��2�n:�T�p����)D��\������ʻ ���&�@���e���l�%�C(�8P?{Da	F8q�!Fb�!s٫6���*������Q�2hl���;�é��acf��a���(���Ԝ��ʜ �L�̻�F����>��!�ܑ�y�%FA�Ѧ��d�zJ2g�.@���BG(�����mp�c@=H=�Z{�p�������h3����X��
�pG�*񏍥�l�}�U��n�s?ֽթoN3�ʹo-ʍe��byf�FԘ��'�C>	�\�9��ؐp����G#�5�5k�7��Tk��*{�G����f+>Pwm@]�"��wT�b6N�2�e-ԩ&�D,��,���X#
������h
s�}�a^vM:�FOߟ�w�6����S\��<O1��xJ#�(!�8�b�����ed�4!���`�n ;��+68�0�"g�bTof��>DEj:�#�-���˓��1!h�>�!p����!�X٘Mq�
�cWD����߭'p�t�Z�W�eDJ^h��a��}�v�üt�����%�<h� ʎ�;{Y�̷�6I1v/���yeh4�+��fZ���-n<;��V��G��'#�{������ܑM�?c^�o��I$ى����%ϔ*��	�u�h��+x��	�D�E�[���[q�:Ej~g�摫O�{�v��5��KdP	N�!��ƴ�J��}uN+��=�#.�#}L�2�t�ZY��5��jz/͠pي%��u��%�8%-XƟ�6t/.��d9�{�z��v�ES(��]m�b
$t0���DY#G������'h�~���|��j�N4ꓧU�}=��[]� ���`6+3���&��X.��xչN�=��c�1���:���?,Z�a�Nv/.k�Y ����i):�Ar[3o��@�JM`�I���C�]�4a1��N�eM7fn�K<Jd?���Q��* �
�U�g�����q�3+�$Mp�h��pc���� �Sc��Z�4�#�@�s�ge�{}�޵Kuz�N�|ܑ��hX�7Ad)��aS�L�+$��y-+h!���,g7eV�0!�ΣR���
�g�BB��u���k����nI^��0��ϕ���}��X��m�Vʖ�jxr1��4ZQ���H�b8��@���'Ͽ���?ш��_�����V�O�N�J@��N��+��24E %����-��/���%�䇗��8A��w۠hȈ��q�}���w׊�74v<��fPdE(�w�3<�K3�J��!���{Oa��2�)~�������!yM$+��������z�� {��W�:��k���(�V�%iS4���Mb �\��hK|F}��:���>�Y�hv�5@_�^�����}��,����@�k��㐒֤��ԏ|��,� ǌ�֛�0��'91W�(n��yP,������:��W"��ɿ�;~�'np(
4�"��:�qSP=��Ǣ,d2��1�\J!�fμ�5�����P7�i~��F�A	V�)��D���%�;t؀�-�P-�4�礌� �9��٣�Уa�i�i�9g��*4�2RzC���r����Y�8�n@�D�cn�V5 c��%@e�~t��J��ݘTu��&��g�>_�Z�D\���_u���a+�:q�T���'��S�*�_߁H� �Ê��9�d��+�߆&��l����G�F3����P�z�u}n7����C�����a'^��bc��"�6�ë��(��m��/I����|{��L���ަDy��I��^D}.[�ʳ��"��³���θ�ԧ�0������QxNT�',�QĻz��n'��6��i|m������V#AL�3A�P<?�*���gl�f����ٸ#�#&�����T��sc��ɥ�c��Q൤!\����y`.I��g!�'��m?��R�%P�4���fa�k�>�.��|�V�����+�K�A��M{�N�LW�7FQI8^)Њͩ�;��E&�׵ 
�Qc:����@�s��9 �s5��3�z�B�(�/=b6R!�P�rGǝC���F_ ��l��p�d�oC��*�lX�whh
1GOU�Ö�v����6���"R�eZ�hr�sG��J]@�`#����C{O�W��V�:� I�����ѓicL�͹���X��&�v�0��=7&�$�L�;����Y5,spWE�n�/������[�,�߯��c��p��d
׉gY�o?&�3�H��X�Ip,�����a[�|�,�7t-���U_5n:`b�L�����OQ������:�{�w$�Z�qAs�LCY�@���E�²Ej�U��6+nA+_�1!���p*�o� m���'�p��?#�1��n�u-�xw�~kʺ������w�2.�ԍ�i��\��$MS�H귗�`�nlC������C�R��K��2�	�b��W�p`�*�Vk���r(f����c���r��KDay���
۞-0dw�ʓ3�YA�/����t�b��&~�f����\y�t�h��b�m:4����4P�ݨ8r :�}�����pƏ�I��na�q�α
��?��|���|x���@�J��';l���������F&���.����ֿ�y�1����o|4K_��uX�|E/ 7�!yDt����x`�24�I����z�Io�qR��l��Z��Te�ࣜ�B��I>5u��Z��&��+
�Uu�M�j��z�{%	�6�j�F*H�Z[��<[������$�_�R�Q���f��_�����S�F���_�52"����3D�4BA5��a.��<I��"Ӟ�3L_�r�x����x���4E`�x?��?�b`�s��c�O䛫�o����R��������G�j�RUp�ʿ0 �J�'2Q�q�}Y��'V23̀������K�lb=��aRi��Β�� �|�=![1���Q��. �(<���a�ɀ��������sTB�y��y&����_��k}sY�KT��\_|�V�p��Q?RͲd�4��쓟D�S�jj~(J3��^��@��#%�Y�s��?����i��`4���6Sq�S��8ؚ'[�t֠�]?#}	jK�v�q��)�6T59_Ϡ�
q��L�"	n�+��܊'[��m[d�*L�ՃS��~]əz��>��4+��4�G�5�kb�L��" ~����$��QŮ�`g�H��ux-_�i$Ax�p�ق�� |�����tYpX"� �si����~k��HS*��u��3K��l
RXY���ʣ@���S����	)͋�@�ns�o+\U���U���԰.P���	�9!��ٞ��/Y1!�Q9꯬G7�'��iL-R����0�
"c��x��6y�(�����3�[�Z9�C�V�V�j�s�C��߅�Ӧ+�����5䄒��rC��+6�@���[R�J_.��y�9n�m�n�Ѿ:��t��� �d�L���3xk��|51�
'^���~��"JK�|�8�y[����0�|d�~]]�o����H�N�{�!l1�kꓺ�D�N��,!�a3� �f�`n>�bntP���p�w)Y�wuW�:X{���#�ʁ���E?M�p�П;6-X��d��*���sO��+ހ�X��OOE5"`��D�h�vK�����p�W=���ߵ�����j����������&;���1����rU���T`��Q[>j�CB���)�H��4������$���,�gW�]n|���R�ؾ�������Phvy���7>�?��Xi��x:K��q��e����ޠ|w��M��0�@�wMڪ��p\�P�ٙ�8x� �#��ʇAKٙ�*�B�
,_�6wj��O�����9b�%���p�n�5�Eʌ�,�w�hxkY�����yd�
I9�x��kvH0�!�O�1؜(�?c�x�s�D�)z�R��m����P���vG�g~^�G,�`k�������ƶ˃&���[����`]�&oVI�=��Z�������Z�6�y�k�2�7x6���9`oŪ}���#F�&%5�����H'�TH8B��H�׌�J!���g
�O=���9�6�i��*M���ר�}c7�Q����Đ��px��4#�3�c?��t��Z6Qr�gz{!�!W`�a��AS��#DH;T"�;-	'��c�s�q���|�s�ה�Ҩ�M�+iX�gk��KoF֚X��J?�*\F�d�|�I��G�Jw*?_RVy�����n�k�0�
��d��yUͶ��-����pz�j�%8f1���1C��n����滋W>�XM���8������~7\�wa`��'k����/��ݩ5����3
�n��t1|Ƒ�(!F�#@�>��
2ǎ��7!(kZ�dN1��hl�4�5~�݂�}��{�W�JHA%�@yÇL�n�%�2�I��,��Pp���i�Y��,ʾ���K��62�H�l���@%qc	���5qe�ޢT,ط�^�����,�Kt��J��R��`cl��� _���<s��q�oe�	j�����:��>Ɇ��-D�,��V��/������u��q]u��_.��m���z��?9�O�q�6��NHN�@�R�
^U��.Z�$2,�y5|�G��	�i�P*�}��+�^P��\�Z��*�,|=�궇�95��ts��=Lo�r���J)�u�w
���7��<�:���"��MV��;���(c��7��2fPP洽���q�<��k�6���,u����/n��7�ߤ�ck������
�������+�L�:Κ�£�1�S�*��ɑ��fks2z�� 5��܈d��Εt�<���$��s /�ʊi~=�9�m�c����&|*���^�#)���x ˜]��5J��Qm����R?v�!vm���p�`� ��1��峩�I�ЫYʾ��C���)�eۉ1��jݺ�肧���#����`��[��[�9aʨ}FU����%���.� �zz�NxtB�����#C(��̤!�6��Jt�]r���3a��5��<���������5�y��A���Eә�pӬ��x�,XHC3�nB�Pn��?��S�))�� ��"��H����n�{��S�x�j��2}+jkr�]����5���#1�
�;�Ç����~\��!��~�[�����V�ٸc������e*�Sy��fh;(r8㜡�����b�I �k��5d{QLM�
�z�����͙�ȷnαe�ӆ�F���ˆ��ܟ᫪��X��,O� ����V��X�2?�:���
/FmxG�"#���=����'bf�TZ�t�k�v4DB���/����; �̝s?/еH�;:��Ͳ4u�F����p����,Ѓ^�v�͘v	P��U'i
��$�Y�f=�����g.i�θ��>����W��@Zt�F`߫T�x1��l?q3���1��0�����4r0�AB�qm<���*!ߊ�H�7�c�Rwf�B�I�L?Fqh��q#��[���6�*�>����E?��"R����M�'�j��Ƚ����@.D�f���Otu�}t�|'|��������2Z1�~��]w~�{�_�pi�V�i&����>�K5]��R0�fWxD�g�ą�Wm�YA�.@�0�˺�H(��Cr��6,������ os��!�	5Q�k�M�)S�`J�4��!}	�_A�ڴD=�;��gkns���Cpf��v��I����R�4f`�W��O�f��o�Z��=�5����8�fa(�H�.�&i�آA��,�;	\��JP�%���֦�tS�6"�k��f��uʸ>�2����֜Pc��q/�� ������@�6��+JN]~F�F�M�~r9+�����uK��uUbIr��m�O��K�0���]��)����5���ԓo�~E��w��ǵj�:u$\���,��j���G��;��;�-ɓ��r���膼]��#1�9��U΃k�sY����:��9���c��3��_�^��E��10��УH5�g6��I���1=�%�2A��"
L�	컟L�b��v-(�yk�cm�Τ��+�[���I�-B��2Daw��䡏� j{l�@e�����V*��ȴ�f��E��8)b�e٨m�\ԡs�P�^��*8]��hu$M�����lf#
��+n�8mZ�0�"�y�R*��{�t��M:n@��i�+LpPTy>�AQXM;��y�dk�0:��r�����d3L��+U�T�)�ᎂu�炚Y��RE[YD� �v?r|��(/'��T�5��$���¿݀��Rif���Α�I�˵�
>MZ��SZ��5)�6��U\L8�19m�����/��5���T�;YV�˦��7Hkk�hm���+ �>�{H��%�o� 6M�蓫�#��fi_(������۱)�
�V������_�ųIf\6�.xߖ���Fb��?T\~�8��Գ(��p�;�t�j�\�����&��$u���>���d�'�
�B� �����"�-���K�f�+n�bBdkG��ȥ��I���|�=4�0#�z6.�b7w��� �$���t�[��M�ġLǽA�{��O�ٷf <PgiO���B-G�7�Ji�3��ssɯ�~%��-�A��*IU2J��*��@�#	�&��S�R�L���K�o�t,h���i��{�@$ʸ?Z|
�\&w1�z�K�����Q҇#o5���':�N��_f��还���?:o��pvj�$��՚�5�Y�O����P�s�5��~��p�^]����>O���spgm����t�x?~��/L�����C���h�׶:
i����>Шu ��Ū�;��%�>����j%��)�J�EpD@����kL���?>%�G�fMڮcK��KrZ��`��D �_������DO��LTy�� �=���u�;B��ȟ�.�t��~����$3�yQh����n��;�K����y�̩J`��	��S�\%���\��X��p� D�c��􎕾�����.m�n�&�E��2� ]|��+�h�r3.#�� Lpy"G�JK|,��6�V�R̫� @�A��X���9֋EHLF�ou.���IT?�5=��i1b��!3q|Z�S����}#rs�:i��*�Y���&��C�t��l��	��IE�J3Ip�,��Z�P��m{�:�#���,61"�_��A
S���
�\Pʥ9�]MMF����*�q�Ǌ��x�;ˡ:��@IPW�[�zp��V���ϼ��Q���+z��'C7\w��<�xf��w�?FiiH��ǋ=��/ �|R�61��L���Aa,NY^	pL^\o�N���!��tUѻD	?vgY�Om��\��sW�!{4`���W�l�8rv�(�n����70��A��~ϼ@s|��frk~"�q�ߴ��YM�i�R������}Gt�����0L��v
3N ����:��
�Eb��>�2)�Z�:��X�_ar��Ȼ7�2Q��y� e|(�s��1]+yT���@���XP�"�VJ��=��\��0�_�É��{������\k��K��9#��
a�#�[�[�
��e���!�]�9&��4z+�S�/�Ó��x]'9g�V�E�l��	�%�������H3ɂ�xG�ˢ��p�������h&����Wno^�Q�0� `O�F_�S�A�)�:et�N\�ߎ?im*�g�L�]a|�F&����ZsH�KE4A�	[��2*"�c��$�2�Hb��e� ,r
��F�>�D��7���a����aS��vQ�@��w���L�o@�@�^���ѣ�{�8����5׆X��Z�SJ�Bk5h{m`�LN������[h�����|�i�D�I��{�ߍ��k�j�Q�.P��~5���p��3�/�6��T���%oTv]��֨����u�v.�(z�쭞�����+�E5�X͝�ʷ5T+i_$��'�
:�?T�rL�d!���O��Ϳ��Lrm�G��ژ�v�ض�^��>�~�@F�8baaʅI��DP n֫�`2��` �v����3J�b�����p\�⌢�ӳ�^7gqS��@v3RLuY����/�-��,�@0�t~hXH�C�t>yi=I�q�q�T��7C�?1��
#Љ�f��L�iak�	���%#���gI½TU$��Lˁ�b�J���|��L�~��A*��������XuA���>�kC������Xf�Gs`���j[�sC���6�(g�vU���w-�L��K!oU��j���8 �$"��_7)L�r�1�A\Y�@5I�xO��8uR?��ӵ�Zm�v�`��5�D�7ј��6�B��������#�g���x��}����Z��$J��QqgGI
+�!^<��Y�c�Y��k�@�ִU	.�y�J�d_7;sN�}/ &�WHt]���Z��$�	���t>*\�����|3gb�oUJX���"x|)8'�)Mu*��+ 2��6�௳A�TڠP>KMc�~B�;{;�����5����B�Hs>���Uy����/��6d�;k��ݤn�(�~�Z�G{�<tu1l�M<C�@W�C�] w�d׿f�%����b'�f{[����D�bĿ���A�_3+iga�RK�L1Tw0n�AF=��4t�����dr��+���d�-"IL����#�//��U���Z�ȴ_��b�O����e��m7����Ov�Wn����)/�b�c�����^l?q�*g�j��E�]�(A�Ɩ�N����Tl�d�Tub��1�������}"����ٗf���Hͺ��<�&?hL7^D�D�o��,I�ʪ��tٶ��tmȦ��>?��yx����4n�H�.�I�ͭs�;�˯��(Q�3������?;']�|C�\�E�r��M3k�3�5(=�TkB0U0���$�7��6�+���� ���P�Ļ΋}�7W΋�4�N�:�֟{�.���v�3Aj�S�YxK��Sw�] �M�`�j{�I��3�����Ե#z�~�[j�1�hv��Y6x��4�m���k�7���N�͂Ҳ�ب���H�RV4��f�g���i�0�(��(3�Wݲ�c�S'�RVh@Zȉ��v�l,kcNm~l(�T��\�Ho�i�Yx��Lz��}�h`��S)ѧ����d�Ďl�ğ;ub���>�*�����c`8
L�JwO����[�[��=�w԰�"��k�:��%ons��8T�QhՑ[�^H�g��R��
p�Vݨ{�~�����S�E0��O~g2+��'�2C�2�o?w�BM�{Vf4�"��}���sRn��fڂ���c�@5��t�=a�ʁ�`����|�F7�t>|_������rDZ&��sB���]k��v��gG
�HZ#x��j"/��@�㍷�|��6?�����Ze�S�"�[
~*HB��d�-�g`z�����bW���Xm�vN,@��og�[�� jfe����Qַ-Fw���B��Hh��_�E���*��A��Q��B� !���a!�(7�{�l��Җ�����μ#QyI�R���1F�I"�Ig�l+��^K�̇ߤ~Z�e�� lt|��#)MՑ5/qV�����\u*���v��� �͇�Y��ѳ�C�k�O4�p�����y��2W���,!�l�8�Mm/L�y�L��W�C�R"M��;��1fm�<�E��
R�2�̴�d�E�X��M�-���oE���+`��+�����h��^��/���F��:>�'�/�8Y��}�:���VT�2�8dP���K0�	])Ez��[��A��)y�� 8�bN���N�N�Xƃ{�=hwC:��l���1X,
�D 酄�*:-A�����}g^@�Dr�V�r�-�*
�k���>4:�tpQE���"��a���*�Z4k��B��nᚪ_0�eV������@�0������vp"ɋ�	���)Y����~�x��ʋA�PH���3^C����9��5��!H�<�x�8�Gi^�5�T���]�w��p����=?��Bn��k{��9��D��i4�q|��"߭��� y�b$N�ϭ���%D�(3���f��y�Yy�{�H(ɀ|~M�_��<�ф�����s;��
;1�\xZ�O{ߐRt�.l�ߐN� CT��MB��f`e�����\9ӨK{X�O���`)�����H� ��p�q�d:N�U�<_cE��c����h-�2qu�5�jv����>��~��S��hh�_�U��4t3@�������yR���%���8��x�ض���vfx4ё��u�_~�.��t�u�<P �r_�@?�~�Hҙ�3�N�y<�Ν5�;�U(u���{�T��iۼNẼI$��<�Ŝ�I��<���V4���^��[�I`�IѪ�6�J�{�9t�xzY�j�|�ҙ��n�x�"�y������� �S��W�Sd�6%Dip�{@S-!���v��(��\WɁk�O��X(����_�Y�ۆ�x^�D���m��m��>z�K��m�����gw�����p��!9|-S�~�b}��hS��y%�Qk�i�����n���������)ٺ�<g�Y�� i�����DL,c�z�P�	R��^Rj$r�@b���2��S(��%x�⟛ڕrY��L���QqQ5�7jh4��
;��c*oo���	����n�> ڍ�����K���֨M���#I	�Ņ&���#_

[Kkh����x��ك:������M��Gh,�rBU�m��֦Ϊ�3㬉�$�V.�s)�jU�Q��Gt�:�߰������tFtW"5��ÄY�����.�i��>A��#�oʉ+j��ƶd�`=䒁nc�@v]�Ȱ�Ч�J�fg��Y��N����Z4Z���F��."������팾�h�▦"�%/!��ᤁm@H�]����R�z��i8�%��]���������p1?a���x�[��n܅͙Ԅ�j���d"|��[#!D=�Hݒ�:��_��L���ΠU���%���.��"��SxM����!O"��FB�Lz��b���B�_m�^��5S�r(�����݅ '0�H��%��Lm9uY�������j����J�Q�xc�*q��>��ɛ�� E�u����kRvc_����R8E�&�I�?g�!%�{�_�gLQf�O�pi������щ�c/O�D<�f������"�Ѯ Z2�"� ����U{�q1D�j���Za��$SSF�x7|�HP�9��u��x\��M�;���Զ���s�^�(�� _�:��$A�ą��ȏ7���t  ��^��U�O�ZB��'	=���D.���=�5	�d�b�(�����	��Mv�,���$
��\7���N�IN�҆��"���Ɠ�im�8}t \�0;����F��JZM��˧ �-�D�	��{zO���e>��5���QҡĪ�����X�~��V�aB�l�k��0�@�6M($G�X2�5� �H��4k#l,I�����̊i�FfL�.ꄍʬ�Z����p"f�~VG%5��S��#��y՗��.�M�Ζa�MnK����' ����<�wűz��3O���/%��u/ŘZn�
�RA�V�U��i��Ob,����?��W(� ��yV`P��ky3$���F���K�Q"�Q�~ ˁ���(1�P\u]PXA�Ɖ\�H��ĽO.�����j�E宭.��ߙb��F'��P�BݻE�.Y	�>�C��b�+��E?��6��=/
�a�H޻
�������x��Hr�Ȓ�lC�1z9��\��R9��5���)j@~���X�Vx75R�o��$��G��g�$��s }�K�L�5ar]65���j�~�����^n�6���|�	su���	� Dxe$N�Ht v{~@�Eq�*�4�$*Ogk��V|M�~La��'f����a���UC���G���r��Υ6�ʩ�0��F<`[^BZ�<�g�A��t���L�NA�r�K��{o!���%3!��Ypc��dbhك���m`��O�c�>CE􍅥�n��.ܓ^��g��
}�4ICSl�>yM�����"o�E�kUl��8nc�m�U�h�� ����q���_�!���rI�ZL�ЙS�^x�CB��2u�����V|��l[>~�ɸ�|�
N���!�-V�šg��oG����}F�Z6{-���W��'V�%�}zc�5>~ _���R)vo$?|�c�����Y�p��g���=J�܆�3�.f��W���^[Z�1l��ں}>$�L^|av���.��](_/���H�# pʃz�,�G��DjA���iX���A�	���d�y�}"׼ �{��y�U=�j9c(k���k���ԇ�
#B�@����>�-����t��"i���8ws�\N�ܹL��Dٓw�N21�ь���f���P��76���Q�siW��*���(��u�>�o���dk���f�ҙVW��R'k�T��H���J�I����jnq]��7���b0~���k��y� m��9�����8/#m)���|50��ՐY�Ʃ��� J��/����e�i�pu����Z�>���C�`>�R�c�RZ�N�C�����m��yٶ�-OL%o��]�_~���m����H%��S�o=(����a��O��i��*�zm��'���A�F���O�wW�=�_�|j�01O��C�GE�����}������s����U���ɑL�n
T�tG�� ��e��g�S%V����\�mz�2\-����I�'���������@%ܐ���E���kN��`�����(:��v�e���V��9(�I5n����{�'����]1F<�#�1Y&onK��^>�.,C7!��)�F�b`�D�m�Q-�	A�)����<�_~�l��6�6��OcϞ��[�������~%��ܘ=�w�M���ɿ����q�|�Ӣ�� ����ː���'x�ט���GW���S}��`]blJX��?�����-�>�~��kO`ޘ��̺�GA�j~H���|�ցⓉ���������&zfp�p2�K';಺9v�7b H}CHeh*f��5���L����'�+I�6���C7�	�#��4&`����T�dcOOY1� K"U�_-���گ�-�f3�Ģ
V���0�a���B�V���g����}'0��ע+�7���=5��o���Szc�[β��Y̥�,�cc겝��զ/�	���nv��zE��ڷ2��F:���lG5���$�6l�	��]AAWQ�+���<��n}hfG�hAb���������	�c�v2H�w�.��ߘ\\Ԙ�+�2wvWړPR����Yb�~ۚ���@5\q�Z��Z�4�3�Ll��J�s2�<���u�9�GB��s�GO��4R����r���mio���i>%�P�u��)�*8���^5Q� �N����j����W^�ǥa��Jp��~��ecB���P�x���t1�e[����R�\d��L	���K��!���c��?�ҵ�ҧ}��$}�Ҙw�毇s�;o�͞�!J-~��-Qb��]��G;E����t��ׁVI�=W<�]��+����,��_B�Mz,�V��C�m�(�OpܪR	,�G�.�sțcl�IDl��5��������ꣃnT�A��(�@"[	���`�����_Q��i���'ZVS��>Y��A������15^��բ9�COa�3bN�! �G3l3��; ��y��{�Ŵ�!��a�Ǆ.�C'��4�F!��B��O*�������7�[���7 w�+c  1�c��]��jZR���䏙W޾��w��~��3{�H����묔Cھ&�n��N�笕6�U��xF�'�W�|�\7T�s��S���ly�
��"�i �� #��E���ȅe�t�Mk�fW�}׃?E�W�&��ul������P�(E�l�d�t#��[��n@r}��vuk#�n�%��l鰑������9zhW�*�`�+j����Z��Ej��J?%�Dd��,5�5:֖���}��ǥ�i-��*
:ҕL�GJ��r�.Ts����*_��7VR|���ぜ��a0���6�'k瑼�F��=馸���9� ����a΂����=ӊ>�
W6�SQO�w��i��]�YP@x��6�n��iDBeE��p�SK�?���cU��ty1�vy4:y0b��H
hrΧr�&VG{
�ooR�g����"�A���#��p��J���l�U�â�7��F":c*P�![���>�8B��@����r=`W�{!W�(��:|j��Q�~�-iơ07(4���i�����S���Wdi��ړ���N7�"����V��௧Z�@��,^�^��r�_�r�i�pvWr�*U.3�r6^�aG����(����$�D��9�b��Q�3_�����"OW8L\��)������s�*�� �lc<��y��g�dZf1�=;m���T{���_ۺ�V(���.6y7i��o��u��Wc�p�spΫ�O�Z���L�������E]a�]sL�e�Q"�b|��3}�|t�3�j)�5�U���1��J;�Z۟j��}��?}4��m���q�q��-�_"'�%z�h����]�n�&�(�\���3��\耤[��ߥN#ҁ���/�<��G�<dxU���>�:W���@m�^'��i���T�9�:ޑ�"F�h��7d�+m�`q��|zw��BH@�`�I2x+�cN����`��a�b��w�y���	y*��r!ꅐXޛ��(��\���)��m�y�д�jo%��Kd������͡��G^�����\�$�@2@�����:ڟAG��"]&��9��EΧ����q6��0*}i�k�)~@�z��z8~��>$���Ṛ@"�����
G3?�\>��[�l�v��%%������Tf�c2��8��Q1���Y���t0�g��w���^i�k0���KZ�E&afUa�,A�Q�~����(�m4kP��s!O�nͺ*��!.QNǿ�4��{@�0"����X�>�2�>G�|��"A*�n��ya�@�xo}C�v��P�R�Jm���f�İ�t�[���0L�����>�5��h�a�ݺ�4x��[	Z�򗠟��ビ˛k�9:�F������8 ��~9RՆC)QF���A�s{:K�;�iۑ�����뢋�$s��Ⱥ��F]A���@e��EX��h��Ob��o�h太r��j��*ct�gv���3�+�Ma�8J�3^D��eK���M>p�rW¥���ݮɵ��3;��}����KGmw���J�������F�x�n���du^�|= ��kw�s�"�a���c�������1��,|�9S�ΛHK9y{`,¿1�����J(�P�vA��UxB\����d[Us�}q�W�.+��g����J�,:��nT�ft�[�)��N
�j�kˁw�шQ:��%*���{��[b�����F$�;�/�U�XRGX�~f��������rd�b��F@�$�,K��Xfi�n^pHV�Hj������F���-
�8�,��4�ɲz�H��jWO_G�-j��Z�����#u�L�5�/vu���P,����R��k�5��#�vk0��vb�
�b�.�q�C#��M��h�-���ODp�M�Ļ�'���GI�i���ńpp��m���_GT\����Y R���NBe��_��ȕ_i"�M|�,�G�r�6��q���ؕ���UGXf_~��d����>Tʜ�w{gv�����a�0&�O�}2�?ꗑ )F$�+X�.���o���>>P-,�~N�>��.k�v���*�q��m�V�@��%�D�~�t��՘l,l �#��P�^f��l�M���,��f\�)�e4@�E����]-{h��*���@	��6cZ��c:�t�� \_���S�ugB?�� xֆaW����%'�{�B}o���z����L�ʙU�6�|I+�ׄ�h^����Ǜ]nO��)�݌[��W��:CnN���b��#��L@]�3j�IMJ��&R��	?C3�DV�<B_y�H�fg؟�YRw�}&ǯ_X��B*��ι�KS	��˅��n�fI�l�:>8s�)b���
�=���6�'�c(�>�Pqe`ҧ��w�;5Fs�c{�%or|H�',9ҡ�l��R������1��yM�X� !�Jk�]���n�^�!n�	��{?]d);_7��Ա�m���S�l"r+p����ļ����K7O�<�=��g��J|N�Z^�����ܕr�b�����a����,I~�����I�,��F51^�[t�1�I&0��Z,ԗ,�2�6G��P�W"�4Os���HSt��M{�q	4���+Q���b^��Mj\�c�pC,���R0wF���a�z����t d��|�q^i �s��7[�qc>�$(
��)u�U���4�#bLJ�֕|�M�,����שD���)���z�;��MP����b�.��w���ҝ*�̄8-�Z�ia�0F��!q�e$_��{>�S+^|Enb%*�9��X-ɧ�ҿ��g���{��&���<��=W�oN��d/:�//D 5�����wbU��v���Z�̭�l�#����j��T��r�|��ϰ\�3��{ޝ�b���vZ��`�(c�;�[{���1���g�e��z("��ESF�27g������[X̋��>��gN+���f���ğ��K�B@!���4gt�ZGl�>�ؒ���iq&է�J�r<�ۡ���Vy�����dub@�&t<)s7�VrQ7 V�鏼3v8Q��];%D1zp��9����'��%:l[�c;�WN
K��n߇��Mt�4[���c��[[�oĥјu0_#�i�Tl�	�ie�f-��0}XQjH�.y ���]��T%Y�Ŀ>g>q�}�.\(�*��)L��h����2X�.U�u�\����w���(�Y/�_@���W�x���V�h��Q^�։�w�;z;��q�-t!u���n��)��3���7���@:����!m��$�۱8�"���%�c)![nFa�y?-��~6A-ZX�g RU������1�F��0�bCkY���k�S������
.q��[���^SA���p)�{^�x|d�-MԞ�� q�.�R���8��8�k�!J��<�V�߸��F�A�K�#�}zce�E�:.���qD���+@����V�x�4`�F�,mc��f"Ԣ*�P��{q*��thw�(��v��8��]��pg�@U=��Y���T�Զ	����ːg�e��hic,d�'(��p�� �`�@k�`M�5ɶ�Q饢�Ο���yx��j�eC��4(a�i�YFa}f���b�O21g�[��qq��5'T8oh�*0&��)R��~D��>Z[�Z�v&M���7�>گ1�[l�K�*��ƛ<�ӦP"����;w	�;5Q�_ɸho���E��6�B2�������P�t��$�[���we*6{&Y���7�$r��^.]E%٩I����X6=Ґ���:謜��"�������6(��<���\�7	5��Q�� oK��1���@���{���A�[�*����x���	��16E �th��^o�-w��:��0�^~ 
J�	nr�
��Wq���M%b���u�5@��^��q`�K;����\K��u��6�jv'��;��h����ڴ�UYD�D�ڱ��| �H�G\H?�ǅ�V�w��˅�4#����^�mCR�A�j��
XX6�A*��G`��t���(�Ԅ�q|���������Q���ۉ��2(�e��)�g�%�@q�Yư�,�,����.�cA�/_8�]�'��H��JOǵ������v:\X���y_X_�aS�&p�G׊2ҵ�!�V�|���U�\uԔ�Wb��0�_A|_��:�l����mܹ4��+X��B�f�L����f��G�+��,zG����Q�'/�+����k�HH�1��o]���x��p ��}�TW��n8JcS[XB��rO6?����[����G�E��5U_��`��3]?�mS�"aK90M���r��7q��@�]�V��tL��+��|�����s=.�{&�g�$�[Ֆzf�jL�gX �~�ԻDE�fi��ܞ+k�2&�f��n(J26��	a7O]V�P��P�a$?8�HAf��\a�$9��,���w[iq��s���pS���G���R�g�����6�E)�Bci��\��U�"�b�����D���z~�Լ@Ʈ�&:BS�Y�����H�K�ȋ�82H 0���r�66)	�.��qAY��f�T��H��hA�L�cA�m��������"!��K�A�.Y����y�8j��8��o<U�3˩QJjx�l� k��-�x7[:���(����E���ޏ�L�|5A|ؾ����T*t�u����!t^}G*��a���Ś��k�LH�r�(�l$p���^ˀC\r5E�j��"��hCɁ�\�Ԅ04,��NU�<Y��G\��c�', (&�-L������q���u����i�Me�8���b6�&��ga����Qn �v0�|�"b��h�cc(\�*'�s�i��^��B���ⶕG���>`����ɘ*���"c�=���Agu#}�`�b�^�E���%G-�{�	Bp��>��v�D�Gp�s�IC�yLd�?��ScYRw<]�,�����H;TB�ҽ\����㈙�(Y��ns�_��e9	�9*��G֫�N[���q�<Q�Sb|G9�܊��j
��=�u�  .lp�5�կI*_��=&9��u�{S�.$���R������;�H�AV�Z�S�AP�:� �Д��M���>;L�����^��[!��~�)M��i=w$��N�Or����D���,�T�_UCc&=���80�*m �:�q#������[y�~ߟJw�H'	�O�X`��O^�,t��41�&�K;]�rF�ף���+:�®�T�i���M��js�J�n튘���#R���4���p�ל���'e[�m��VE}{��G��:����6�z���j+:I�b�P��y�{ɿ�<>~�y#Y�ңK�]0J��j�/�O`މ�2;I��_z��3E̡�d��!�m�`C��is�1C��o��"�g�=y��՗�J��qf���A��::���/B@�/7o}���ၑ 2R)� �;�r�ha�cb&gӞ�i��.�\��~e6D�,|W	��M��
�W���'�gq�P���u��/Ҽw����(.����6V�O�����0�&zY=��[���ߏ;`q} �©��!�$�?*��Q����>Bd��+^i Gf��Ւ��C~���qP�ٓ�۸y$���;z C�B��MO�����@e�D��{ֳ����,�t=o���6'�}��{G�O	�I ��T绌��&��ۘi���xϻS�:�pq-��&�~���4m)^x^�L8���t�J�ŭDo��#%�����J�;e����xi�T5J���}����%0gW(�$��oV)'�=�XcP���N�D�B�6�b����h"��8��ĥ�v)F�s�����k���]�v\5���>Ѳ�q�>�<�I�Vxt���.�E�Bc�*ZZNV���4.HH)��C^���Y#��I��ħѝ
�P��1%;?h}�|tj�߉O"* ���qT��!͂9���b����$�
������P�M1���KslƬ H�|Ah��A�k{�9'��>;ނ������`[ʁĚ�:jDxO��-;� �2�e�ɰ>H���j����&�qa�z{� ?r�V2�C@|��f��� ���hD���=v�J�pNY�)���A�	�ZV�8��~}92sz�/�²���`(I�b�@Ii�;I!N'���S����gܢD}�m����$�÷����w�CgO���垑'�2:~�t���fd�7������օ��[�k�u3J��}m� ����ٚs2�݋[�t+��[b�̦և%J� }7�#��>ji�y��.@�̀�o)+ν=�&� �n�@nmj����!:T61�s*�$�|"'IQ@G���ǜ}ĩ����Z����b����=�S.x�?����S��]��2�v���긲}�k�JVk�$����d�M��G�-�'����T>�N�d��&��"��_	U�S��L��Ր�Y�c��u�!�abC�š�D^����?����/�iG�8D4�@n��u�7���B� �Q��?�6;���,��k90t��[�TC�:�4��;%����{�XȈ:�>�����.�Q�B��m��J���T&��r�y���,�ؔ�%ά�b�4�!V�e���l(^%?0ً��߂9}�'$hKaa��l��Q��i��S[�HM���꺲�N��~�x"�����i_a���'Bx(������Ks��w,;ٻ��#�C=極���o[{�B��
i�����+D����R���)� z%�λ���: �f��(D�.�I0�S�8�8:u��T���!�O�Y�Mhv�'���<�W�`��b�q����bD�ʴ|�=Id�B	nC�=U�i�:�"�Q�|!��%]:��i�8%Fe��8���c�� ��i�X���-���h�ݵ�@�PS�+�I`"��T�n�I	�~k3�����6�j�4\C@�in�w>�co�Q'S�`��"��o���V�lp% ��:����l��jdo���MA!��$��ο"2�w�t�2��t��&�!�~�g�R���1���G����_��1�,#hq~WX~�%�;�x팚5�Κ�-�i��.�#�h��y�#����Q���Z����S�z�s����cH��Y�>�UOM<����D�v����t�t�/s���F�0g,��[��������=��8�;̴��&d���;�y����&�Y��QV�&���W�IK����?c�q���~�C �|�y�7��ѕ�PƗS�U�sW���S���B������8����]�7P$�'��#� n��C���i9�?�>!�ys�N���3M���9WU���]'�9��V��']%U)S�~��`mK,q�gf�Ʋ���v���7ѝދ�L��(��W�fE~}�P��Z
��?՛UE�\�跜�5˿��k����KkY;L��B�-�������	hFR��e���\ebg�(N�Őhw�nn�;�u��2v�%0
���0�������g��@�ݪ3#F9�~]���.�f�N�1��`�����mW<��Hh�ϴ��o/�ؐ�w�6)�r�N��[��d���h�S	�՘��1�r@��j"�#�l�&�l���ԭ��f��5�k8Ͼ�`��>!�^�(�J2�20�Ƶ�tlZ�w.r��-�H�H)�z*���3�SV�2�fR����c��62ѤE�8���l��E�|�]��#�Ӗ+1Nu���#7�R@��6�v��P�}��$e�ǻ�������2�7$s��ڴ��7��. ���y�Fc�`�g���x�����u;F�[Z��ZH�+�B�w?�c�	f��+���	�H�Z�:h���I�2����,�#��V���_�:1�J|�|2��}��{'����o�Lz_l�����.aY�����v�`�}X�����Kr}"�p�z������~���������;�l�/��{��$�n��H�-^zL���'4�"|W����Q<�V�M&G��-M��c	4%�2����+<n}�L�B��!�r��h�̓i��Ly_��Z��Zd��7��@�ʘc�i�>=W�faxFt1Ǻ��gaw�{ܚ@ƾ���g�}���84��+��K���-h��G%�n���i9j�"NI�T�^f9�m��֘���"Pv�Io��~��hN x��^4�d/sB��X��Ů?#�9ɖ�����G�i����n��d�}<5�M��j;\�����]�FE�j2'JQ�ǩ�e��dJ`�V~��X��dSt+=4�ɡ�Tl4���=��(�����ў��Ґo�GC���Y1�[9�FBjo��୲?�@2K�'�~���s(�R��Fp)�ۊ�UX71��s*��fj4�n �W̞ۤ�䏭7\o��[�m�`I��L���m���H��^�h������2��3�k���������nو&1%�>ӹ\9vT��U�����S�(qL��_T�\r��6j/8m���b��C��Q��w�{6�iu�PyX��nfZ���0���
�6��K�ؐ�G9
�f��\��#�6}�O9R!��j�HC��|"��EI���?Zz{c���D��~;j tyK=��ew�0y�B8_+	s6�g�`C�������s��#���o
jgS`�@q�+��<Y�V�G4���3`�kޘ3rwdK��±R�*I@���"˂�
>@?z �m�t�m"MY@Z��,[�y�I�`�	R�`%JQ�������6YR�YF6�!_؛=�P�bu^h�bu���EKK^ؓ�.��5Y8�#.�kP}Q�E�Qjܿ�ʷ��vڎ�X�m��i{��H6���׺jJv0ӻ���Gt_�z,]�Dr���Y���c-@���9��3B�aY�ZxU}Ռ f����B���x��
�z[��MdͧB��`Q�=�^Ct�a)Ƽ�G��j9��i7?V+['�n�gb���f�b?n�5�����s��vE�λe׾JP��1�3����	ۡ}^��5a�ކ��=�3t�� ���d��:轘$� �$�����2�#jke�:b��b����:�3mX��L
4)�UZ��g�<�1�&�%�6�e;�-��s�m��@����H���&u$��s�Ȱ�s�L�!��R�w�hz���P�7�h_4!K�ѨsH�E������㡺����sM($ȱ��|TnGu��d7����$c@͞�N6�U��]6�٪�qa6�.5�9����6?������~56����W��)*��5��`Z���� �J�Q���c_�)�qPZZɃ�-�z�Ƈ�g��Ȋ��4����r險e����[�{�����Xˬ�(?�Q"�-��jm�6A�Շ�#&����w{�����5���6~�N�rPC��4 a�q��t��0��S�z]�0�?q�r\'���-
)�lB�,�?F��4���-�(?�:���������^����]��,������	Z|�"Q��6��X��}�����X��Jx��(����Z�T�cĽ���s)f�|$#@�1��}�d�o�Qݥc�}ԝU��1v!B�h�sT��qT>��c��n�r�}�����$J8�0�2���xل��7�&6O��O���}5�,��#)c�L�@*Z��g��u�m!�[@��]7�����4��V�f�E�������*�����(�����Jۉ��@̽G��}N�}��.e*+����6*��W�Ph|��T�T���-*��c���/��`�=�X�!C9�z��MT�J��1��-�\e�"��6[bw�����z�Q��&8̌h���1{r����:��(w�I/�/�� K0w��7����&!��t��$d��%x�y1�I���[�.':m'�B���������)����!���jv��zg���V�ċ@-^��-� �)���+�P\U��z����݉� |�*�!KOn�{	A�X��}p�v�;�����
����?�<\R]��[��l(6U��y�y�g�X��#��4V���������l����إĆ-�C#A�~�wD���?�Zx�Ӧi�6�5�/��
"�QC�+��8mbE�W�yM�qR���C� i���K<L�]"c���|fR���F�u6n���\l�EP۞����*#θ|{��<�X����
 ������;;�X�âO��j�9����������~�H�@���~4����oj�I  O҉X�j>��YP]�&�B��7�n�*�Pa!���?����.q�1҂]��<������Zb��=�q�{�=7�6:�ů�c�T/��^�P�����>Za�((K��������%�f��i+��ڹ*w̎%��9���@�f=�P�����i��<���`O����Iȓ�Z`��t�SA���W����]?�n���K)��;�h}W�����E�⦑r!nV�d�Z���V��y��U�=Ph�A3�����D�4Ķ���z�@��vQ���y;@Pϼ���rY�-�&�fA���`��@�K쩻����j7Ա�O�h�c�䍟�VT��U�݋�|$<wc�0첌M���h�^"c�d9{��>-�0�!�:�ە�͡*�C2(V��m�ڣ�x��]|9vdHh����G��gw�����:Av��ځ\Rܘ�9(&�^�41zV-状Y��!��O��}�̗���:2
�G�#�I?<W6},$�McK[]n)��g��Ĉ7�|?�m��z��jx�X�Y�h�9�Y���&�G�h�X���b�pA��TV�b�&�Ja0�i��o�v/���E�b?4�"����D���HY�ԫ�)���k��<*�c����f��YStQ�W�ʉQ=k���!Z �4f��t�ē�UPVw��;������*qʡ'z����)tG�ȃ�^�I6B�˦�U������^������C�@�kP�S�y}�T���b`�����o5�1�W��w�E��	-7�|%�AKO�I��F��n��m�X�w�wS�Hn���K
�POe�]Eo�NyԾ��TS�X��>�I6 ��t}!^���2���K޺z?��Զ6��7�!�{���ʕm3�x���6�+r�V���XX厴͹\%���d���/�0v���@�N��oW|;�(m�����ZM��Zΰ��4=�1��-cE�=Z���cY��vJ���1*i�0��q7'���U�F���c��uWC�� @�����[�AW�'C~� ���|�O�1(>�,�m :�{	��|62���+�$����1��Gn�r��;�ߚ��ğ��t�ҟ9"1`8���ӽ@�M]�kP[�A�2X9�����u`i�a��$`dIPxż7.��Ts4V5)9~�Væ6��T�j����K;����	
Q�^€�)U�*C�l�s�u�V���.��ژft,n-�k�N��l�C�0�wG��,Gݔf6�Ћ�E��\c�[}��B69Mr���<Vj���9hcU���)ώ��4�&���J��|��m({!@��r���������t�j�����lX$B�K�> p���<�q��Ş�{A�S���0n�����	^�4�)�2E����@�ٗ����Ӂ��=��S%7Z05Mvn +T �,~��}P�\��� �����3���$���D�Ꝑ؉y����Y������b/jrp0"�+s�I؆��;���1."2'�&F���o��A�C5կL!vT���������*�TP����%r@�~�N�L�t���m[,ke�� Ҭ�os$&Ie�Q�m;C�lEÐ��
0��,O�����5;kdh�-es�@�
��p�kϿ�w@e
8\�nͅ�}�)P_9��8r�h��3�O$������YZ���2v��� N���"�7��1Goc6�l�,�ռ���P�M #����������֣�#�����CZ�:p�̺9�g�1�i)���`��'8�7G��8V���^�z��S�-O�!����Ķ�?���S��ٛR�?��=���k9��׻�)�Z�voJ$�w:�q+|!��H���f{�`gI��mI��p��^-��Э^r���u�6A��i&<��� �j�B�yC�m�o�%	N_�b�r(��Y�Re�u���N�k�Cð #?P�P��0�j�:)����ǅ��A���X-�)���;7�� %��'I-���7Y&��ŏ�3�v�����!�%�wvY�7}��DO��E�-l`tx@�)��俯+^6����_�˱_��o����� �ۥ3�Y�i�A��B��1ӿ�pB�)%:����Ƙ���:KU2M�w��Ě�*9��!���擬[HR��L��t%��Ol�wI������S%��䭭�rq��#�����rq���s)� ��|�5yx�zz�	h�7KklaOyKK��C��q^�h���"�=4���3�g�4��Q�9�T�6�RRn5#�mH
E$��f%a�J+��L/��'�Jۺ��n�;�Z�~ ]�I5���yH�����S�S��N����������⼢m�-PN�DT�j:6�-G{��pC�ɯ��L��DY��o4�ތf��#ïWV��<3��-��x|��J#�\)f�ь���x��<�h��H=�x����I>�T�`G���3h�TU�@�c�jE"/8]c�K��Ia4��{4�.�x'�7�%��2~�V�q�<�S��Xd-,�b<f�s(k��UF�ꑇ�:iYE�h�jwA�T�{V�\�ډ���
=����� ���U ��Pi����Z#9��&�/P��Sn8�"E8q O��Qo�DW��/��?��[+��!��F����M�a�8d�){�C����!%��S��*JF���+swj�	>�SmS�]���_+�?1 &X-��Ȃr�	�mά��/ց����\����9�2�_XDw��'r�9>Z���ѪN�%�u���|d�ޝr��>_��}ّS�`�qvPZӊ��~����<<#���0�`;[hP���V�И�K-�Asz�+�߭�tL�P��h_A��uCr�3IM�i���CC?��d<�bY�H7+<��@����MFM�̛ccC�_���r&�?��\��E$�At���`EX@��B�n飯�R���hG���%׷$�h�M�R��,��=>n�p�rN�W��s�R�x�U�Ni�J�)�c."ANi��ъL
Eu�I��I,�%)[x��c+��Ѿm�������)���Q3G��*��G�����(g'�?S�WDro�::�۟8V�S�n�O�]yMںͻ'���B����zZ��G�j�L�#�HEY;{�����	Y�Ƣ��w1N�:�"�|Ԅ{~��/���Xt����Nf��/k)�9{���s�����O?YB�\a ���{�����&�epUz%C
-��dJ�8[ʻ�3����B�A,���� �þH˽L=�>[� R�9g���M?g~��UV���f�y3Z%0f��H>\?.��5K��s��L�'$��8�Dw����_�����6��� 5C���<0��������X��p�0Sk�Qo���ʦ�u]�ɲ7�P=K�Qn]-�b�8�a�arWV����֩+t������b���Ɵe��K���@�J�O +6eQI.M�"p�"�tRS:(UMv���:�-�lC1�g�b�]��t�,I���@���R�_1�!W��j�����F���9�ř����ߊw���X4�>��j*�X�c_�����k�A�[����xI%
����ڲ5�z��I�
��t�lͫ���7:&�1�X+1s"7�����.V��'��n�z���Oj�2��WD�)�i���»nҥ�o���U�j�� wQ=�*'���P<?D���v$�W�{K��"g%zG��.�W����� ݐ�&83հ"5�F��A��Q����n�!�B54Q.u�$�V����D��mcdK���d�D�	ǌ�V�@���-��H*�t�� JM��!��M��X�[�����{��^W�x��}��,�)��*�o�	v\-en��[�à
�)ǭ$%^|׋s6kyK����9�����K�����/���M&o+aԟ��n���zwiюJ�"$C��h�/�����\'_�$�q��9D�`FM"�����NX	�v[�t�w-�J>����頏�uAY��8d�n�|�	�S��5ǯ��D'��<�3j���0<���b��w}��vzOl:\ޤ/��?}I,�����.��:�$�]�wX����>�u
dƟ&6��)�W�
��0������ʩi��T�O�h��dD:�{\곔1��v�����`��O�������Q3��6]����k� �ͅ����U��(�&a#��Xj�|�!��Ӑ�jf��jj�*]��1�յ��K�Ԩ�4�j���:1e�s�A1��D�|��b��}� ��d�;܀_�x�:��K��kA����L3}�u_��c�y�MM^�(Z[?'݋3�juv�I���I�z6[[����L�`6�pi)(7��3���a�m�!P�dQ ӟ�+`�IB�4��l���#��=B5/�=���}���
#lK��(N YY�M��a���?L�m'��:��ʷ����2h�O�=-/�E�.C��mYBx�'��sb��o�'�]p6�xdjF���_�(�$��يt؈����FK3琫�K$�������/R�|p�TS}�2�aRo���ђ~�xj'[�}[��2lN!.�b������FN���~�Y6s�.޹�>�u(�(Ne��gn�rΩ"��O�r�s-u(��R��þM�u� ,KH#|�,�LF ���]�������C�D�D�)s�.��'�+U�2?R�HO(g�r�D��Y�6L�[��"���j6ҫIP�ܭ�҄W�)	�d*���
2�?K�G���	��B-��҈k]�\��D>�#�\�p�sz7��,��V5�&�U<]��������x�M�c'5�gJ�p�x��^<�B���~��|���	L̦�!�Y�鄞���e�Z�qѧgbio��"��ܘ��h���Z����.*Q��"Ul��nl�����_~���1 ���ԯ������fŏ5�LZ��@h�g�JI3 p���
4}��kO7�qȁ�t��;�z��~��Q:2�W*|����Q�,'�9B�u`��R���H]s�ڥ�$��ɾ��)�/ ����spdKP��M
p�:X��-�K���-x�R��G>��;�n+}�����s���QW�#�??.�oA�\*�s�P�Q����&�j��M4�{�b�A7��i9h���#���RD������Y�ݼ�NRXG�ymW��5J>���a��p޿d"D%�������wW]��5B�JyC�d�v,_ێk��h*�l�俚Ag`��A�8:�"���Y�c�P+,w�B|ԓ��:�@LUS�6��W��0~��˄�\/F,Ь!c�� ������$�,�|	Cu�I�[=A��9�<��3d��Rh#���2�O� �p�������_F|�S�S|I��������0
� �&A +�v��Jy�m��\Na�`��`1����rI�uƮ9�r��(�VJ}�&�ԧ���]�[�S�����ј��H���0��G�������Gz@#�D�u��� 
}x�� _nHS(�����{���l��c��s�@�\�z�j��t�Q�7�i��:lyk.N�1f�:�0�WD/� fכ|O��M�F���Z�ip ��1[7���;kləfH���R��(�(ǯH�+~|$�����M�ou 7�L�⃔��s�Z�N̿�hNE�W�qƼ��`�hN�t��Yd�(Z#��M ����;|XO�BQ{ܺ����]N�M&.:��%\,
�P�q>y��rk�- ��x��1��\��@�p���gq"Y���N���T
��z$R�B���H�zkej��ʶ��b�/�����G���fz_e6��-'!��4�$��N�!��yf��4#񉪶�M�S-[�+��4��uɬ��(�}(`%��	��UA�b� �$Ci���'�����L��ƊS�J�5�429=�DF�ܪ6r�NZлܟ����ܻw�Nk��}4�v?�141ӻ<�v���zw,@�5�n��a3�w�~���P�g��i{�*�بy�a�f�
t)ד�M��M	���e�	��53�����:3���ኁh��<~]$����?��F ��i��Q�U�H�y��i��3 !:��ѩ\Am~�,��߽'����'���5�Fw�sEn?�S׶�Ƈ�t��B���&��l<���z�A��{�0��4�a��p��"[�Cپm�]^���}s++q<CoC:��t�� ��;���a6�Y�������d��nP}C!��&��IPzUxv����I�`!�Y���J멅�=����
K����1d��Vt���J��ݽ�@jY����=�4�R��)I2Bkk�	~�݅o�[Ux��n/bR^�fi��+� ��)g���o�K�����!�T����#}�����ZRU�/��{�5Ky>�ܿ:�m�NԈ�u�D)NF��n�!/��ڹ�ca,}���zv��I`ӏt�;D�f«���a�m��V2�\}�r �l lYK_$F������VhH�?ů�!|< ���_J�s��}6�+`*���(�<X�i9��I˒��fM/��!@g]�3����:�lA;:���((�j� �ϸ<�%6Y�u���	�B?�P�L�"�w�w�����J��Q�5`��3�~�$@n�W팫]Nm�0<Z--���1H�lL��P����dmʽ7�m���N�x¶��>VX����V�\������m��ۮ=���4�����g,1]�b\�҆���Kfa�46�W���eq���l�����A=K�s�Dk���m�I}άH8�}ǆ��X�ޚ�9�{���괾�B��%�tn�"�����f�ϻ�G�����5(3��9��&�n)����@6�\d�
���گ��>�I#�tCn��rr���P*��<S&���&���n�J�u���X��E�t�Qn��2bO�ϵ4��ȭ͒r���\�5Kf��Y�f@�S�VZ�4zEk���	k�zc� J���M�P쯩HN���ܳ[a��	�V��ed��-�2p��%��+�x�x��I���Rd�\�2�ԧƼ��d��}����	ĭR�T�!�D��|QZdA���' N�Gl�
��O�T5�O�v�N	�독MV�Θ�߿;v`����-K]��2�@n���e��}?��fra���9阚�8�Me�CC�-
�Ы�)��.	�v<�rwhD,�J��7Hy�6>	�#ч��o�rvm�) ���.&���ǦK
{-���L��#@/��G�o�[�:�V�v��.��(��틣խb�&T�4i1*�U"����$�geK䨑��=���W��;I�b�Yn��#Ԉ����Q���t���5��@���H[��Q"�?�ى+j�mczx,f^h*?��`�Y��?tx0���N�ƶN��	�}����b�dЊKl��=hz���7c�B@�$,��X(���K`��eX���x;e��c×Ҏ�ˈ�FJ�	qf�}-�M��(���M�=�C&���Bp����׿&��Ǫq\�>@Z����F�����$z�Z<2���q��]r<R���#�j�I7�N&�R
}ä��(��������eW¼�n���Z|ǶQ�?3���3d����e >T7�|�/�`�!r��Cĭ��A7�M��z��U�` ���u�t��W;I�^�����PL[X�n%���G�z,F�@T�hD�`L��P��iE�W����g&"-�L�3?��9���ԕ��p�P_4uZ�a��۷n"���3\/J�{����X�U#)�֞`EQl]&�Ȑ)p���hD�ځK'}2�(:�
?�]S�W)��Z��:���3�<o1Л�!I�U���- U�ۂ�?W�E�D�ڻ�ɴYJ:�˶\=9To�����]�G�xhT�2�b��x:���
���rx2�����;�ވ��	Ё�0>��F����O�vMW��<ۻԣ�;w���YE+�\�O���cú��lxV5K��C���3���5����N�en���7�3������X�`f����L��C����w���Q1:;�ӂж溳ܑ���t���߁��a�����7�ӭ1U��'�J���َE$��?�;�@>���eP�ZŊqRu��^�'�N�Y��`�2��Jrs*�sT��h��1�Rw!����&�BsL���ܔ�̭�s�,�^E�{�y���mh3�F�Y""���ai;M/i�S��N�a��:�b�� j��O7�� �)�D-x&̸�q���W�i�p��ǥv�hakkEh�&�a�m�S�������Y�<���{0.: "��S�2�5Lw X1��/p��q�K�����R��Һ�f}i�N.]���jo�0����ՀFv���t
sn�i�"7;8��S64
7��7:�Z�����[854�!�@����.E�x�� �2��A��������h���-s�A �I�S�lc;�(�Y��f��8U�[3f@ՏP�&`hk�Ti����ס&V�  ഄI~%9�@ϕi4���$K�%,n�`@$[E�
��>��R>�ܰ���E�f�R�S��-�+�����P�M���ln.��oh����u�Hѡ0ŧf�x��y�4�����r��X04��q�y�1Xh�����i5{O٩_�� ud�wk��r� ��r2�Ъ�G&JZ f��(x(�qz����
-����]���4�d/ɯh9��NX�*���򪈼��F����A�ߋ������R7av%V�,�/wg5q�f�n7�+Zp�^Zp!0�����鼄Rs��Vw�9T���zX���d%�8�1�7s0�ҏ6Q*���AQ\��� �	f��xʩo���թ�ȗ��@\���J=2YS��K�$.��O�cg��u�/��DyHoVn��Bv�n���n3� �VR��(Y�o���
���&�Ep>7�65ٹ:{����P�Y�χ\���Q���G�X��$(Wc�3X���a;�(��H���rQ�>�Ww<̃ �$��ʅ �C�vr.������������A����·��H'�(}
�N���;�e�P¡�'�٥{+��D����E	➔}j%���\P%d��l&���;���
�N_�#�ƴJ�ߖq�]d���`�^A* �XXڲ+�1�"���n���V�?�jg�����!�|�*[���R�cB��6_��Ҥ��-8��[}�D��6����#��������U���3҅.�:����߮{M���43�+�=׏��J����l�)1��*�C���8Ɗ0��Y�<z�Jga!��q��z�{Ŀ��'���x�K��o=�7�B���4F&��*�x�S���!z�o����~4��F�񈈧q�e��R8<�:q؞�.���<�_<�5�-�fƔJ{�V��������g)� Ft��2�����U��R)�1�Y�a_��p���
�1E��-f��'�5P�b���R�)umA�V}���R���!�k�bOhT�1D��&��X�E��h�m)bވ�V�b�������P��э�h5����o}�N`Q{R�i8m�R1��]5�v�)�(�k`h�WAt1SjUy��%=�w�7a��j7�ma��C��݉��ú=?�Xts��Mt)�2�;Q����Ω>w�����݁�:t���*c�6����� k�x�(ˠ$U/�f���7(�d�15	�f��~M>�^￼s����(#��@�|�1���gY 	�ZGCP?�Zkn�@�tQu��ڃ{�����յ�#+8_7�������,� 
R.��W�����`��'L};���:l�8E3������~�֭.'M�GdzŻ�{��G5�/wn�#f�.?���#$�w2��J�,sH�\�/f�����E���I�͂#_�4�Y��I8n�H-O�j�����*(��MBf?�.�5f�PS3p=X��Q�����njz"x�'��Dz��D"��U�)_d�����6�Av�Ay
�kz~M6w��`t.��)�����q�on�����^e��=��8䂷�Iή��Hz�|����pIf��_Gia�!!sc�s��8���w�f�����'���S��(Y�[E*�x�M��]J��� ���WI��i��qF/��|0)Ff{�XF8DQJ�V6&�d�eu�߰]���^�BMm�ձ���+��I(E�>�{������Ʉ*/�Dq	���`��������x]\�����n����ޠI�s�|1��g?DS��_C��1+·m�<r=LMoAԺ/ ���B��bCMs�[*�B�GW����M)OR�1㌈c�a�y������~�>��g@y�� ��hq�W�M�A��W�O��k���
��]4=�0����!��t2Z
J��B}%:��n� ��V��}3��~�~��i
��y~��b��1���6�M� �p<g�撣7w���=f?d1_���f}\$o�v������P��\Z��>�;�x���⇠�+��<o<I��̂�ʊ�hX�>C��!����!CR�T�+n�9����X�&ҽtz|�������Ե���5��
;���L���M�\pp��6M��r����3Ǫ��J�8?���k VV#r� L=�Dz:��C��µY�`d`�'���Bۼ!��7͔U�d:�e��~�� ��9^5�n��v����E�0�$��.M'J#�n4z�ԛ&[������zhM	�t
���x_���ѩ��T�\,P]�퉬5�#��U��A��+_%��ņb^�؊�e��v��v˾ĳ���b���/�sh�2�wh�����3mP$�����%:m�����Y��*)�χ�q�8��>CK�3\M:��Q�������M0G�2�5[+���w1ߞ�T��O<��xb<���$��vr���_9�J�I���y����=�V�@ML4�l�a�^���"EO����5��G:5�p� �/O��x��v��/�@���+�Y���?��qxs�	�7�m�fr��3�(`�j���$AdR�kS��}S)5�3ݧ\mV�'ܱ�카emt�s����o�DAOpq���{G� ���p�/�D�R[��&�W�4~�P>{Ç�Mη�r6�`�-��n�g=����*k]t��oB�����+�9�0Yցd�Q��(���nK�[,J�g��!��N�@Υ�u�bgv�P�{�*�<c(7�	$��Kj-ORƅ)y=Y@}5�j��/�x��􃍴�:)��gP@�up�uAf��n1\�U�
����K
a"0�R��U73\�%��V�v�U'��o��d=�
`�2�w���ǋ�e񼾃1ۖ�#z�(=Ev0�kT�F���!|2J&7a���R�Q�R�[��e*wA�RE�l���)#���t_�˦�a=�X��Yj�]�fXӹ�[�^<��P�sR$8��e���}!��;S��ѿ����!�T`/��[����k�~�М^b�?E���îL��.(�G� �'tq�`��~ ��x΂�db ������5bpz�9�WcX^�߁Z�w��A�:�^5���J�ة�\?���A�*C�|2¹�Ӂsa��.���9�
6����޲�H���H[������K(��B��͔��"����Q�v��/���������cP�`K��ܟH����[��MPϢ�4�0+?a�[�'X��6�����^�k��)s٘��,��߫ޒV0F�B���)>�����̅�T	��q�|�H�)_���/�	�Vㆻ��K�bG t��8� ٠�\�x��x:�"E3,���g_>A�&;����'������7�v\�-�hn�3~��s,�9\�L�͚��l�|�|���Ͱ������^cq)���x� �Հ7ɫ��a��ޞ<��R���	��@q�Y��w�T'��|�-��`@�=����)����Npt��8�J9
o�8w8����q�*S���ֽ����L/�M�(vT�����_�7�\��`���������ϙ�[�"��m�^�^��H^!�~��<e�w���J�CsӁ�
:?3u�&���X��dt��C?��Y�@��@��C��0�1C�Cp�����Y������z9��k��O�.���ţ�J�������A�����p�x� � ����.�-��P�����U��.6�*9gɯct�����#[=q�d��Ķ�u�XM+@��^[wvf�Ɩ� �!-��?�/��(?Φ �7���NiC2n�u5����|�J7��������e��ʐ���oi�%Am`��6d��9v`�p�d����hz׏,
RW��:�ƈ�J�d5��X��%�������'(|4:��z�����@��Lߋ��$��.�-O��#4�]�o����٣-�Z4�`��d3Oi�MĬ�4��(m;�s�1hF�f�6M��0'�����k�fr ���|Z̃�L�PLͧ�S2��:���9K���eK�XfS��%��ָ*L0ȧ��7a8t>��������Ř�T����2�+��b3�*1K'�N�q?�u����TI��K�������X��4/P��@�\mLv)��c��~@��~��f`�������7��p��ֵ`�������|��5G��,��E�x#+�B�r�ᴼ���vh��a焿���c}D�G����� hLW��hL��K��h��e]w�g�[P7?l��Chܜs��x�����?zb��ܻ����EAӽ��_N3~(�xQ�U�d�|�����`!�P��;�yG�/��;���I�]�aI?I�ggc1k��)�<��ϊ�9�}9�YO��>�&�f}v����z�6��Җ�ZB\��������h^�V,��uʞ"dH�z�861��"o0q2��Ȩx	���+k*}!����p��)z@��B�0����9W:ڴ�m�]�B �����u�1�����9<����w�� ��Ê�������W�@$W8`�m�zTI�R��%�q�[6c�1;�©��BJD2�w�~ѱG�K�b��v4>�<Ҏ��b��@��m��f��I�m����ȝ�ߜ�(A�9�+'���?�;##�>�A�ߗ)�rn�(���^�aJA�ɗC3*<	5��+d/J �al����S�B��|�e�iY����!�Ld}ch��	�r&��<P���}&�2����l������UMj�4gN矼ԴH�t���
�#h�&�f�����i#@�2T���^�.����-�IN�|G%j<�n �5�0a�j��dXk�f����D�m�f��Q=q:�{���X�����%��C�k�>���a�Z��P�FGf]k&��y�}��:�Sz��g}�|T���̟�i5O�t�3�u8�$b�$o�N�C,T'N��.�L���7�=�X�/����mD��S��;�zN9u���ч�}��@��h݆��i��-*Zl��F��oA�,�-k~��qNJ�wQpa#ZgOA��n��٦�s^S��
�Q�pX�Q��
(^�n"%�)����I�g�Ź� ����
q����X����A��*A@��Z�`�*jh���Qa��I��	���2�����S�Q51;���t���"la�Y7��n����e�֛*�5��)�:���_�+��8�����h��kc�3/���x����pkZ+�=�=+�4<׽3;+�|h���.����wY�J�jl�(+���YTԬ�ۮ�4P#"�'����K۰h�ձ�	��t�o�G��e��&��?�>(��V�7k�]h�$����!2.)H�����ţ��Ƭ�����|Y���P�� ���,O�H�a	���%��5����:�-�ڀ�V�J�m���2�^�΅⍯�O������iNş���]���N���T��O�*%�j���0e�<C���:��Y2)��˂�κ��R�*C[p�1-pH��~��^�Z��c�&����b_�TYΈ���+��9��ԍ�NO��&�?�CV+��txu��o�2��q��T�\���(JI"5������gY���0�WS��ͨ��{=�x�m{3��oZ_AS�L$�?9N�S�*�T�j��q�W�NH��)7�|h� �����ɀ6��{�&D�S�G�~F%�!Kpi�Os�Ǣ��?w���d�->��Q�蝨�8C�=a����zcF�����:R�O��k���>I�#��B۞ :�c�k��EX��2,��m7m�!v��A˙_�	����(�c�#�G�ʸp���B�����fO�g�V��;GeF4B�x-7�@3T��(pK��*�����Ȣ���@��g�\[ =E*���ظ��>9�ŧ�:��#���Ĩ���dOK��cb�Z��.�;=,ntz�ļ��z�A����Hr��n�R�H���_�M���?'���;�+~QE>���/�BԟYO��|��C��5j�x��Q���ʢ5h'����a��0�$�7�I�����>�ߴؕ5�&B�xh�雦?�^����X��?��;�Lbq�~����x�
%g�8\�r��`��%���I��B�Gؚ�w�{�ڊ�C�����x���tk�3�'�1\�u���..LɗT�(��w�C�����┖� '����J������a���h��ۣ�Q��8V����Hڑ��N&G��*����|������0¶����t���9�$%�g��?֒��:\3�;��4��a�8���C~�ulr@�=!������#��A��l�)�&`
^@�� s�E*�Yb>�T)��A�SJ�a�	n��jI�B���Z��(-����-�I�Yk}Q�Z����J1�z1�h�9��;Z�Y�3���:v�!	������Q���Jp������c#��� ~s��e��$���J=^�'?$r#��3t~}×�,�Γ6*��}h�f ��x���ra<K_�ߏ#�G��#7�˫4�L
ji�[ju`,�ĄުLi����R-D�6��8��9�.�h��p&a.���!=𢽿߅lo�48��&h;b2c�6�$�D�^�	��GBR�QHW�W�p�c�U�����������\��ʳ�sk�g�|�b!K{a!��ҽ67}�5���S2I����äX�?k�l,-�E`B�ѰM����ρ�;l��M`����F%�Ȥ][�y㗥����3{K-@��rM��>KQ�m���{fŔ�e#$���y���|���`F5<��<�5/����\g����harQݠ\< �(�H��襄h�ZI-���^��Y'ˍ��X��Kb׹�-2�/ b�>�,�v���f�Q��k�o[�|������]M��>���<�.��m�=x�^,��M��nޚ.i��R�. ��wv#�P,Hg��W��J���q��X8����H�C��M<�PS���V��C.��e���x��~��~06ɥ�.-8��R�;��=��A�)�D�|ͣ�l��`V���K�ཽ�VRS�(Y��L!X�z�}�����~�l�,m�bk�U��~�&X��t^�ZQ��c�b��z���L�He��|�꫶�����~�����?���t�}�7�a��B⯱u��8�o�ҧ礖�L|�1J3�rC��vW�e+�0�PY�0�B~�ʵ���>�ʛՇgp$=� ��ͦ(��0Ve�jҳc{nN��j�n�h��(Z�q`��h��hu��؁��Ð����%XI�Az-C�6MRx�[�,�o&��a����9.R��F�����h�$���\�\p�α� iT�d�I����UZg��U����Mxs�n,�,$"��E�����������?��u\F. :+ �/�Q�9�W���(�$�vJ-��o�hD7�F�ZlN��,���F�9�?�P�ڡ
4P��i�*�}�)�LT\e6PdN+�r�{M�7��%[Ҷ��&f���������ݪ�kor��g#��s�R|%�]Y"���D�C�j��.���T�u:p�>tnD]]2xY?eՅ\��ܻ�D]��5��N��^C�%���o	0�q�
aꅔY�\h,��	�L�jWBc#�"���,�"k���O���W��Иy,z�T=\� ������ |?"h|Iܑ���63��W	 I�\�.�׍[���xu����9�?9���+�.S|��B~U9%��u�#��c���v	Аܩ�'��O�VX�Cx@!�~��',�;-�;�ۧ��򀍌�u���<�g ��5�1b@)�"4����m�Pv�[T-t��|:�BBw��n\��we�6i9`uL�;�~��֯�R-,��~�p8��Rs����ѓN��2^�Ƶ;0lD?���@1����vU����晅!էfhy����:�s;h�壨�+��
+�u"�&�Y=�-�]@��K��J���_��������L�����Z��j��1�Ԣ����v�h���V�򨚶9)|rx����e��%D��v��O}(@��x��RYۗ�V��,r��_�h��+�Xt�4�#���`�Tٍ����K3�+'�&a�"tH�Z�t��})C2>�P�	p�~@&h��[�J��p3}�^/�6"�S' �]:�Пrp�r��Y��G#.�t��`��L?6��47O�Dg��t�8�S[cܝFkF�wPW<��N��ߦ��%>n��K��RϺӆt���^Mm}�Z"��ߟVSEp~s���q!�����w��@�~��w��U��7Aa��2%���jRFW(1~-G��' ���-*�wp��G��t�X�eݞ�^�wm@nXE�7��>��g���}��G���l]��x��Yf��mBy��HC05�����\w�c��QB�&DU��
C��٧�*i[.ʑ�F�B���r�*�g�^����e�m��hmv�����"��XX��d��� ��	f�����@�w<E������n���eB�k����C&���#Ϫ��#-2������]��6l��z�&�jL�a �q��R�׌��i+�g��d���`�Di�y���k&ok�����I���+��U�C���Ԛˁ�u��4
��e�����:|�-=s<)M�G*�:����'�� �Ee�6�!����$o����.�ɫ����W�D5Ң��O����7���}�l��F�i��$5G�5��N�{13��5�/K=�^�5[��f��|>�?Nwa����m ˞�M�z�m�ﴖxl�ؐC�.1�n�IG�Z���m���C��K�v���!�x�@y�R/��>b�q���^:r_4 ����Sjd:�k�V�&�<��놙E��uõ[?�[�~��6������N��G�*����Z&�V�� ��?֐��;�b)�6{37�2s0���n�)|���wIy-��~��B�ٳm1����E N�1�9�']��nn�;��|�t;�VW�dϧr�;˨�