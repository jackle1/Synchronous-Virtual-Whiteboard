��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3�[�����Pٵ&�����''�qe�-�?
�%w$�W��[��m�w�xH�O�I�	�@����[oVʭM�A��t��B�gx�K���8C��G#h�̾cZ���8���L1�}�L�RZ��L/��W�p���;lB��*�Y��4�%]�Y�:�b�\Yv_f��!P�{
2G�-�Pi���xhB�ё�&���7`��G%����U�^�9���t�M� ���X3���#���u�鉾μr|Wh��h��Kɟ������cG:��9J>:���ϔ"��nE��2�����>pS4s��	�(G4{(S�L�:U�.@�|R0�L8������j��IB�"���N������ys��ė/,ҊN	q�v�Z��\R�w�0xtʎ5x5�������v�7\M�k���%n;c-<�<;�`.���B1�7���[�D�\�A��fIj�)����懋�f�7��ǟ��Q���eO���}�D�^��Ok#�H��@@�
5KPZ�Lw�<<+�?�^�^�ᝳ�0G���(��/.���`�2����=�2S���O��'���>63:�\��yZ�{���]9�#TXh�cee�Z�VH��ty��Z����8���lA�<����p�@i�ّ��|j���`�1b�N���nV��_���cq+L���6�ݿa�"�ѹ�e�d��g���r��͖��	��cN]l�*��-� ����/��5�?	�D6s�����rB��Co>F���]�&MQ��R��=�tXB_�*\퍭7��������q�^�.���%�.��6��TR�B��L6V�0uW��<��ؽ�<:ن ;��#*��_�_Q��8�LtğՍ'����b�l�u�
LD��l�^;ϖ�]!듓D���)���"j�/ �@&�KGs<T��}�BP)�<�$�4���R{��RV����aVl��ڲ�����p� ��2��z�؃v#>�t0���������`�6��~��ԉ��?���&ϝû�"�z�s�T @N&�C��'�����%�XKA�R�i�B��÷�[�Y]�%��R>��
�v�)	mɯ\�=���p�	�k�ܗv��Ыk�E7�G�D�&s(ͥ\je�c����[�Q�*s>�-2��54l�ܰթ�\�8a��Y����Έ��T��O����F�5al�/�=�p�J�τ���0+��#tK�뿫��*ި�o��hط�O�'	���Iֶ��|Y���a_թ�X�ͭW�	�o�"���8�Q�9[��u�C��/��$
�"H���ԱQ�gw߅�zM�r���g�!(v}�MLb[R������b��R�p̽NA���ݑ���>Os�wL_��h@d�aY����_ʣ�o�!�������B�G3u=��.�ܠ�T� �98z'��T��Ľ�"�M�?ߴ� ��1�'�N�r�f�����%gQ3e���d����	B2�1��y?��X��WSů��m��u�`'Y~��Q��1�G	'�.�p�_�9R�m�$�]�=����L����B�� +@ �]=i.��D,��ZrN�O½�c>�,�NWk���G�|�}ɜx�V���,��B3-�UD�-��8����2CȎ��H�o�6kG	�HI���R��9���oRX�'��q�۽4��%�uS��s�Шl��\��.��*t�T�ҳ��`j�H���H��,:q���I�5����4=����E9<?�<:��x���ʪ����0�|?Qy⊨���O���D�ݱ���V0c6e5Oe{-��jc�W�]�-�	2�
�~�-q�!���U�6��O����֩lL��O�K�5�5�ڶ��N3�`|��,[�*�'� ;��K
���ľ�+�mq1�C�=)��@�YNc��'�4S\��*�l�GAc�|����69��*��٠�'Y��
A( ���I�+d�i��#��P���{�}n�`s�l�ɝ�-����`Y��S\�����v�su�ՂX]-�V����e����Gۤ*�D��؉���55g�A�<�<��oۥ/���c�����;�e��H%i�s�FM��?���,h��Ɲjbt��`~k��R#}�U�o$��(�'��A��6h�1�)HQ?��Wc3�s�����#������|����?��R�@�'��x�j���m	e,͉��ݿJRVթ��x�)2�/ծEքJ�{!�9?����J����U��<B3:)�=��ǝTL�+qn�99=ȑ���;�CA�0[���#���k;���S��Z4V�9��0�2�@��	�v���M^v�a� ��;il *�  c���o�DP5k=[��~��ݹ�g\U)l����Rl!���|N��j�,�@�j`����׽��|B��l0���*����?�����K�ߌ>���PD.������U�qG���C���Qի�>�V ZfT)jl�1:�9��w��/D��{(���` tnl��ĵS���gZ�6����~`��+�L���y75:��� �_�C���c������1����5����؈M��u�.]i�<��a��.��6������ �B���NgL)�D�r��6�"���ږV��2�KIC���GW��x�Ƴ���"æ?�ￍژF#����OMR6/o:�'Y�]�o�_��W~OnI>+k+��c��ݨ��Ȉ�����~�bm��h{����?o��wk�L>�����FCJM=M�W��X,Rs#���i,8�}\�}��=g�R�?
+��Vd�ۉS���]�M�帨U��ņ�L���O�XeN�m@�fy�G�}h6��K�ǚ�c�ݣ��	�6O��N���AOa(��O���[S�y 3E�d�C���#�mU�[�6�O��Qg���m{:�2�U��讆���x�
n3O�+���͛s��~�Ւ >�BH_���Xs@V>��c-�=޲��? �WS�	H�P:(��1���mF[��������{��\���D}�N�@�$�'e;�yF�þ�N\�0[���|���V�?tj�v(�����a��<y�Kf���iΥ-�̓�풎�Q~K�����&u.B�� 
���3�)�<4x"�� �M�^��k�T�uų�	nyn�E�J��l�Я�~c��.�K�pp��̈^���v\;�>ٝ�7:��͓6ʑ��̵��ّ�G;���!X�Gi_ K��1�iIh�ap��t��l���#0鰝�*%���JN���9�f(����]MGk�֩�o�y/�Ҹ5�˕v���*��ua�{����)BX��?�sM��2<��q�X��G �+�==�U���H��l�=1Edg���y��.�ӂ�XR�3�T�t=��~��بci�8h�3C�dI�q{�	9�nJ�����4�n&nM�<[�Ô�b���k=r�&�Ǫ$���z��߬�죳E���)�i��i�,T)�ڊt$Sl~k��Z(+J�⎅A���:�w�����V�\s�A����ϊm��H���y㔃��Q�n6�;=ܩz|5��;u�o3�]m�1{�DO�l�;G����������^�jx���T���.]�X#��M��Zf�dcC����_=�aO�.n��Ɉsha�f����I�+�~��4��Δ�NL���`�~�a7+��lcZ`И���9�~�}�3db�\�!�����l=؃��:��M����l8(`1nR��*E�Y�ܝ�:����)u!�������gc�;�C�1�PzS����^d-����Z�f��E�������9+���4�W��H����{��=$/���jBi�]������c��}�jXaMF�M�F�;n�\O�zX����+x!��A����Ws��{-k@������'t6NP.:[9K�&eQ��l�ZB�&��5Q��~z*B�g���f���-����"�H遱xȒ6����ɁY6��f��X?�e0���K��J�K�f��#�nux|�G�Dhb�ɲ<���V�"��}zPc����}��Q@'@�O��t�C]�T�o�,�p���{!V�ՍqUOn�N3x�:�*e�u��7�i�4J䉞tZ�Jo��W�d:���Y��a�+��!�T��=��w]N�ivzP,�NrO�傮z&�g��)Qs/#4:T�.n~Z��l�x^RZe�K��r��-cG��ë��El�&x�5=@�!�\�M}�5��7�)��;Վ� ~tJ^�����Q�LdC(���s�����(��[%~k#E)1<�҃ ,���,~��/-�X�����gԍ&H�g(��(B��B��m�W�a	��$��b_�;�n��E����� 3Lҳ�V%0�V��r�-3�㏥�O��l=�G�=�s>�\^Qq��KtHX�[!.��&r4�>�H��H��&��?D!�(��������f��tFe�6s��گ�������Ќ�l���e �#?%� 	��[���m�a��H��B�������x���I�/%#yğն�z�qu��2~+��`-�C�C�5��!(���w�J(�>�(�)}j��)��=�j��z�r @��m����6QKR�mN5���TYˍ���j!�[�Y��NR��Z��'��q�K%����o�/�x߸���u�_�9@� ����Ȍk׎J����;h��q4%�դ����*�;�2{VBJ�C^.iWօ4+u*�K}Y�/�WnG�41��S^g�y_=��:5�y��o-Xc�*��$��h��R�+�ơ��
����L�ȑ)z٢�RH��*%g�S�Me��)k��6�!� �3!��@m��JGb��
�j����߲�S���w�K�>���=jh0�}x����i�ڼ^��P鐙��2��i�6���r�?4L����Z�ػ��{=6>�볮=��E�b���l��38����̾�ͳ��G��^�fb�o:+�!-��x��jYQH=��#� ����`C���a���`�Q��Хu�O���p5gh������S��<���c5'مK[� �}�TK���։���VtK��CkM�A��p5E��J��LQ��Ԅ�)���B6���~,kjơ�I����l����N?�j��4�)e�pg�[<��^�B;J&2/����}��An���#���}2x8o���=�[�&ĳ+��F��e1����]����_�5Ksg����ϵ��g�|t�7��m�L�3d��a,�ޮ(�<���(�����wJ,��r���#�����^t� �����aYĈ8�g篸�v�w[!�d㚍�?��,�jYP;&�y����Z�$��mʄ���ɂ���]2�����t@�G)wU7�R�Y(�C��8�A�5=�������p���Q4�h ���2��Jm��;�R8��e=BS\���}�۲T�:e��b�G-QaQ��"ܽ ��& 7��s�t��s�p����ŉ����]�ǹݶ�u/v8�!�앟Ԝ5ʹ��z/ڃ�x��f�7��)x�v ��o�������nHo茁sNH,)(��������i(� t j�����Y�D�@$���d�Y	һ뚌]��p|~�T���X�����r	�毁��_'/�9�	l��x'���gi�?&6[E���@9���(��ڙ�q��6{�VL�w�Ⱥ��%���0$��!���Kz�#ZږY-�H/~p>w�s���hi��_2�(�T���I�����y�нH�A���@�(�w����d?��6KJ�{'N1�,U��l����OZ��v�=>=��D�(򆅖_Bi��cYoٗ�W_�����"�*zw���.�AV��R�P7���t������%>Ό��fG������-OI�ͽ�D�y|��ط
�Ds��f#+]�E�z7o�K$[��r�wJ��W�?�8�z�6[���"XX��	O����4��-@������B/���l��W,NG�їsB�#6��Y[��Z���}�zO�\��FW9��E��[��8i=*Ь����?H�^lL$0V,z���|�������n=T�|��y�7.ʦ�{���pX[x\�k���=���>��pP+ <�.)��eiOơ�(>���7��Z� Z�|��{�ߐl���ӻ�&_�[G&>�[*fX��<�o? y�WB���\��R��螾q&����q?�1��5���kL�����������J��]�`���Yq��b�r�7NՂ�+`( |`(c0r��JRǯx�4����(��o?�+R��Fp!�D��.G�Q�8Oԓ::��y����J���%$~<�� ��H��zb�����5���<����~�l]�S������|���#�>�G�E��*bV�n�E*v^��>�v{��o瓗������eo�mPCr���0Q��&�vR�؝r�(�&�#QN"d��}j[�mF�ZBr��ES7@O��r��A,�2�C���y�Տ8�c���-`cm���@�(�Ќ����X��Ņ�n�3��TI%�����[� V,8�.e�1��j�xMg�
؏�����m���$��sA�Y2����S����`f�Jq�Fy���=�C��qH`R��E�l�;��p%�+G��z����qO��	#IX.���>9�g���`����/"^�6$�,�����ʎ����~[h?�YE˘�}�%��m�t�'�r^VP`0E�ekZ�
���A�F�!T�
/�?,E��@X��;�q3�Lg��������Y�f��wһK�*����	��K�p��  >��X��� � Xp��률��/.p�IR #P=���g)�Ϻ̯(����у/H?��?��O�G� A�:��`�ǫ�'j�R��>��]X�]�SC�g��*d���t~��@�ꕡ�A*���ׅ�C:�q�q�ſtՔ�����{|^��Su�doBf� zHZ�(����H�1��b�m xP��􀔁�'}��V�cA�\��+�?47�������x��l��v�O�����L|��OqE>��Օ|�;��^JP��.j��O�D�#�<�u����t3�Ki������݁�s�T��؍�Һ�� �CL����ZkJ���M(�;n���:�ۮ�g�j�@��U4u�8S|w�����X 48�D�V�\{��zLir��	����#�ԕ�ru�W!t�y�+��Hl��r���j�@I��\�;��b����;�g�t�s8td��<��w״3�o���;��"q��@ n]q�����3	��>����Y�`�T_!���t��us!�� �ϥH�����xE������T��R�V�+�C6�y�Ժ�H2����À;��x�ఓ�AT�/�#fgNP~A�2fwL��Ϊ.����h��GG�tLra�q"��S �S��gH�$��5��_K�!1'Y ���ya��QwK�{�iA�v����2ռ�~����lNU8���04N+���_����	n���9m3�7���[������[�O$�W 8�u _q��D��V4�����5����xq��Z���e�s&|�BKH�W�H�MJN2>����/�V��Q�[n�F�\�Q"�[�T	_�����"�B�e��0-�k��[�n��6MT�[��]u�h��Q���{�9�wę����TS@���O��c")���0cM��e$[�)�XQ����$*�ܘr�� �� ��1�Nv`�@Ǒr����$ܨ���U�v�u�ȶ�ʦ	[T�����&GM�Ϥ!Z�C[�A=��w�E��ҡ&�5�����qQgu+j]&��{�)�Ͽx�]��h1�<_�y�B���{�W���>��x"���d-ה�����H�6V6�:7�r�{@���3����*d���3@���Y�O���>�Md�xUX�H��>�/n��L!4����"r��>Y��d��Y��l/�<( j�{�F0Q��=@u�C�(u��䪩t��q.n�M�3ת@9��s8]��`�ox�T��f�a����o�DU���RJ�WjMR>�	|-����yCw`�cνPt�K�QT���wM�e Ȑ�ļ�׿���6���:x3$g������^K9�{{`D�l�/�LЌ�q��*�N^���vm
(�p�>yd+b m��I�S��Hu1Q·���ZWKj���z?��c_�}I��w�}9M�5�y���B�E�Y�d�H,���W�"o�T!}�ؾI�Y�0y�nw�k�t+q��_+K?��#�p�*2�=3<�GHL�J؎Ԟ �Ȉ0ֈ]�d(I��Z@2�:đK� _�u�p�ଋ"7\yp�ס}!R�C4i���].����%�rr������tt�j�GӇ���M�C��&�eo�������ƺ��G��"�[%��3.ʖ01[��񇉦(���zn�d76��Q��]����=	���m
A���7�������ର�?3]����Mz�,�Un;���R��@�����PR�Ԣ������m�����٬F�C�3 }4`>!M�d�IZ`E��QU���N7�G�bo�sg��AX��>����OQŞU���H�gb�N,� ��س�lwu�Y9;�Υ)���\)T�+�׶|������.\�LM��v����N�,K5�5#)9��{�p�gN��
�lÌ�RФ�a��h����e�s�v�Tl��|��r�
[�lCd��[l���6�c:�;T��h3�f��ŬIrF��,&aƍX��h�`�}:_M��0�p��H��35��`�������Ѕ�R';=3ɸ�s`��d4�fLb��E�&�U�&�r�/�s�qɛoƓZTտ� �I�0 �>`�򇫆z����6��d����f�|����DY�Ԥ ���[�Q1G�X%��+��y��F ]*�J3�ףF�U3�$d���
�$S~.0�Y��=$�V�wjrjQ�@cK��W�3�2�����T}����A�^�l�$H�'/�t�{%[o�	#r����θ����`��ɑ�>%��z)�$�|d���TI�7F3���课.Bh��`�l(�m�2& f%����.h�5�1�HL-[~~�QU�}�&!7P�ʻߐ*[C�j\�����VV��ۚ���˰�E���/�+�H�ǭV�J���|�Q`S�����_4:�R���5�{��"},A�r�>$�8Q��Y �E�"<�����i��~>`�>��m�H�VA|PW^gpP��9!�&9�x��1jȂ�޿"�*08�"���tP��� 趠k�@�9u"�z���c(��?�A����	����qߔu�	±�+�ԁ7�)�Av�x�_K2�dP��(b�Fp��rU^_AzLv�Ж�7�K`E>�w�Ŷ��\��B�Pt4�9��i���u.U#(��d�K������y�__&^M3��ߦ`I�$�CQ]7��%���?�^T�o�o|d�8�F��	I��A;8�������;"�w��z�+�#��짂�;�iH�Sj=IS�Go���ݢ�DK}�c<Wg�JWl�/M������t�tBICy�^�WN	���(�tM���o%�h�X3O��xf)}i�z�Ɯ���ͧ���-���LJ�Y��1��n]7l������W ��9o��~����W��$��ל�� [S�?Pe��9L�g��=�z�L��N�l;��e�}�uZC�(v�1�s�&s��EP
п�T���s���tK��hu+�d�~^����u�5{O©g���=�aҽ�w��p�U��ڇ�׼��&�Y�| s�E��Wb� h����GGN2���.8�x�K-�&��&M��4#SD5��9�hپ��Q�l~*��#�
Ǫ���B;���N&�!�9"�YxA���g�2%��	��H�"B/m����x�4��b���]_/b)?;C�#���dS~����t"?b/nFϪ6j����+�LK�c�+�"����G7e�r�a��ܒ��i�����c"Q&͚����5ג?X|v�_�H��X����g�?R�^�l�gDճuR7#��Z�Z2-T�Q�t?�2�:�w+���~�DQHkl�A�;��X4-2���PLzs�qQ��P�^�c�f!<VR�fN��]ӈAQ���vp�9y��Wܢ�= VL�\W���0T�֫\�q����S�&ɿ�xgӇLȲ�[�(���R����E�޵>�":��񯚦+��#@�} h�p,�OwJ$�-7�t�N{�h��	��>k��+|����Qj�b��i�'���w��P;� .xư���ʹH�/K��Tf�G�	��x��&��z1��	5_]%D"�!�H��,��Xh#���.�j�"��^ֈ�me�cn�u0��ڗ
�^K�~ r�`����)c��kB�$�_Edౡ�\^��,�QM)a��!V��v�v�eۍ����RR�F�x2�B*d�VZ�Eޒ���N���mB��f����*�M���/�#	�I;�:�����Tp�x�i��1�����^���_2�>%v��0O|�E��6qOFXJ�\���Z{Y{���R"� �4G�4+�w��K�i:
0p�|D8���D�������NJq�F���iۓͻIG�P�����ZV�2d�+�c�cQ�<��o������J��k�_=v�0��@}�4�Alטp�&b��G�T~��ʂ�}�꬚�H��^�=ZZf�hQ�w�2���e.�[���U>>F���9�#~�\c|����������(�%�3�����-��]��H�'�V�f�}��+�0�MϮ�js3}���\������6���Ȣ-R��+�X֧FnB*���`%��W]�T�$^����0*�������'��2��v�.
'�6�+�'��`�:MTl����B������+H�t��8��F���"��<��/��'�m����+C��FDjr��C�5h�k�|o��Ō��/����穿U�6\
�>i������D59 @S(��R��3s'�0� ��DMc
�yҬOco� 뒓��ReO薨Sͽ"��¹O���'(����{��,g�hI�<�
��.X��tM�.ʱ�x�;_e��V�m�,>��ƆF@�<[7�e�F�J1͎7[c��\x)�*����{�q%�����>��2-MD�C������S�J�l��+�Μ1^���^Օ�N�k����U�� 0��+��`:̳�$wocJ?*M�pl��ԥ�װ�b�;�WLӨOC}�ʪ�P�W��'Oݝ�6[��!���e??�$��p]L��rb�ز��1�M]��iֻ8;s)K����h��[ʘlhh~`PNW2���O`
��S�:N�̣Px��
,���{?`��t���}E-;u�t(v	$��\0��.����{SM�&E�3���|Z[�C0c��Ƶo�p:��w9���ch�?�h����b�Oέ}��t������(-����NW����Hc-s3��e�8:'�d��\�P<-����7��>��C��P�$(7r���ٍ�2�(\M>1���S�-� ���S�2� ช�s�g�N؎�U��VY	�u���N�Sh�I���PgY�ĭ�N�������i��Yp��U�R��	;��1P�i�s4��wةq�F^KXňr�o��bL��2}L��j��;����@��l��BVgVfץ��x&���=c��5v7'a[�f�"I)��{z:J�0Fr/`���<Ir3��y0�~��-�ީ��Qm1<�I6�s�ʪn�E�𡂚��� ^B�L�a�[Ra^ao���D;�Mo� �@8���
���L�xn�fg�����Ѣ,GF;��\�GuhW���|�]'��E�B���!F45[ʗ�n�P�8����5G5��Cz�rw�V�=Wq��A�S�d����ޟWY��B!�����T��֐�L�5����ch����-�h.P�>�eh���cW�fC��+�M�+!�����Z�c������g�`N؋������.�ڟd[\6ۢ��u���[1���u7�2,�0̂k���Y�}�k�kP��;��)G����C��s7�k���&�&(N���Xj����X�@�Usa�Ed�J��B˺�i�u����өޑ�tZ_J4x�� �����踣k�}\]'9�8 )a�-|󘅈N��uT�+<ޣ�T��*a3����U%�"����n����C2!�����m� ���b%Ahp+�.Z׼�<F��Z�@L�=}�Ԗ�R�<T�X6��f��Ne���T{����t�AT4��p��#g�z���p����Z�lS�+����r�j|��܀�1�H�7@<�ϕ��O��d�k7W�e�Tk�"�C�/�X@zo*xx��U6���̊+5J�i�$�#�$��Ng#{Y��c�'6�$9A&Kj�k�}+�e���4r5���oPӛh�v���~�B"�؛�t"lO	�KY+�	�]�QϲM�b|��-/�2"��Ћ����:5�͞�A~��p�-�'�P��_q��'�� ��W,�}g��=�f�^7fV�=@H{��r����%���-f�♐Α93[$�I�F��L���еQ��Б��AĥCB2}��5��������r =��Y����5��Hc���O�\�e�/�<��\b��NJ�'��z��g���D؏����,J+a����)q6��2q8��B��'[W4k�������9E�������u�!8"�NTi~�1������%�H���`a�F�#XK˫PD�/)'�h��MR�{ԅt�d:�he�� ���Boq4a�*���s$���s��sj�Z��	�IR�ľ8�A�Y�c�	�a%f���Z��1�@��&����,��v�)�D�;���;w�#J`�2�d��p���>6n��M�]3��t��E���&��ڃ<��
���{�El���ʔgٟ'�U�
G5LQ�x�IU�f��.G�eOi���"-�}��f��|�릉P(��<\2/�
��Z����cqO����u;�#G]l���5�h���D5�OꖴU��A�5�q���e�,���F
0Q��ִ=�����!ɊDFO)��L����y��)>�&:8R�h�����<aזVVf��NN$���Bo�;��'dZ�H>k���9�NC2|������:���'�jQ��:�����%� �L_�	έb>�T��=��DHM��7��~5<f���L�+��.I.�e�	�����o�Hz�����Wq�ҩv�S���*��\=:�/��������R%�bJ�C�����)�0�i3D8E��+��U�I˿�a�g��$BB���~��I�a#c6`�1�|�C�,���hh�\@�uc@N���2�k��*� �$��1$���;�L�狤�s�5S_V��>->�
P���v���v�׽��s�ļ�ك����B2$x��:g��c�P�Vԩc��O�tu��d�O13��=�n�
�M����ί(��Q��s
�c���np���t~�ߔ���&�w�Q/�7!Y�l�/�T%�����S�,���	���RV(60K���,M�"c��]�2���;�UY#��R̊qU'�tX~Z�Nv�W)���幁c _�,�#�܌B��㸵��`AZ?�,F �h_��#�ck�{{aR�o���� V�c���0��dWx�)y��ʰz=�m��D�7����-�:�;�)��7u]s�`�%Υ�q���s�
�q/#�+%)�BVO���0)N��J�v������;��Npg���E��*�K��{����6�e]����9DiEt�V\���+�� ��cb�n߈.g5�PDzs2)����x�_��傳��S$��\�X&�&�?�v��C�A#�p*��<�U	����۟��=��O�`Hk�*q�S��Sf�/�!��Ӽ%�@����'q+��g� �o��P@(�����#	�zs�}ج䜬\�wMI
�&��ٸ����g�j��H�gM�G �V�z-���n�:�}������r1O`G�0֣,��8%��~��ZC��,6��>��r\�c�lLǃ����@T{�>����S��C�<.�!��Y�;��j��R���(@���X�=�u4�S���+��K��E��z���@G�TZ�j �	ڧ����LC���H�2��
[N�t���L3=�O��@4�K�Zi�9�iZ������_. A���%�N�Cv�T�!�*��k���\��Հ�bH���t��Rz�,)	�N&�y(<��Ym�,O?\���M�"2�A����e��Y�F�^a�����n��<����q��0��r/�<;5}S��=�5k"�"I�A��sT�T���e��ͅvW��"�˴��5I���U
�4Lx��G�@6,W��J���BӬ�;E�t��������S�t�Hi^_��s?��F�Ae����u�O���#cE'������]m��3��%���=ox��,\Ö{�lz�ϟ#���D阜sm"�d�@}o�3���х�!r'���ų����`^��u_�q�q_�j���vV�/��:��A��nN��0�O�y�A���&Y	�[!�4t�j���9]�i:��`�����H��*TK��ED	tP���A�FD��Lڽ2e��������Ê���W�N�h3��&�i{�V�99Nl��E�����L��9)�j��'b�R� �d�fw���)R��!����4����=5bE����i2E,p ��1S��w�M��]@�R����ݡ�S�Q���Z�1�CeT1��-=�B�,ZDp��6�Xh_`���4l�W�Ə������"�}���QRZ��5qbx]s��[��A~ )�덶��{|<��G���u�Z�����9i_s��&�RJ��`:`�j8bpe6�t��;�g��~�=�QM�I�sq(ɒ�xg��fF���r��c��}���;~��]Xn�˲�C���)H��r�,��DI۱B�
�����g�H��L+����D\`	�2R�d���sJ{.+ @ɞ��_ˉ
g,&O�tPr�@o�`��x��v��W��{����$B��i��d!�$�(&�1�S�#�e�Sî%f�#_��c�����H��(l�{ş��E��2����BX�%�pkrw����jZa2d�v&���Ta��'�eE�X{8�w:���C�kg�ټ�r�1��]z�$"�;QV�aU�^j6#	�u.�W	�Z�L�*r��iWC��6�(�m��q��Ѷl-�����%��2��+���!}1/xk�MU�;E=��g2c��W	�������gYW���v��S�H�;�8���0,N�O|0��blo
{@5yenz���[`.�n��5�xt�۲�`����Q�o]��аbcg�8��xݷ@�La@Q+0�b�w]T?bU��I[Iuq��qYH"\����-��g��eD�X�7i���RSD�)���a�)#:��W�)��
��_3����ߓ'ө�vi���7��C�@n���}��d�ޠ���/�S`N��(�b�\Y�4I�v[*{y��5X�>gv��p�Lx�q^;�A�Ӈ!{��j,�Gs:��6l棍��|\�q��n�����J������k�F,��E	0�����>y�އ���4���h�pu�� [,��#N!���!D���ā>3�B�qz�N����Q����>�y�]�Nj�Ɗ�..�c�li-�BoG���Q�{���9H�@-3c�9J�1H>gGI�#�ٕ��Iv�ڝ�~�K
MŬ[Q����*�nH0��ܩ��w��D:�����^��O�S�x���u������u���W���9T��ۜk!��@�� ���yܔk�o:��B��yA�m���|p���� r�8b���7�v�i�R�+)���@M�k�ͫ��럻��e�H��ꛋmN�3�ʴ�o�V$	7dbB��������'� �L��'W�HKx����߹�F��O� �[��U����Ч!�9�o�F�QH:��� �<�[``��!�F8(4Gb�q~9�iţm0d �/2>'��[��6��}�0J5���L����W�)Mr�����7i8˪���4�$69�7Dyt'l� >˲���ji���9�T��;A�v��Bǩ�ga'9$`�k
Ѫ���1<?ɹ���j[^")��MF�fK �n��X�4�r�w��e���N��,�c/�@'�|��*����ߓ7>��/A��ѷ"
В1�*�)F.aZ�-K�������r�K6ofR�{qgB�[�}e��
hfnw�DV�o뽫�b���q,�
��q�/2�KK\'��`}�!K��s����e���(8>��J����R'���D�cc*c�+Z��XH����W�Z�e�h�?{16B?���;K6K�]�ܳSv+�ף���=�x�B���(-�G��}Y_��R,��A�����[���С���G�򑺨u��}~@�l�M��)t����+9�&3�KcTţ�y����H�J+���6��uD���z����1�d��YV��� �����@�,3�n�8or��0��g��̥� �X�\,@F��,�������s�*	p`wW}k,��S����8��L���I�k"��;�=�]֖K.��+�����dP�����}'Mq}�rR8�*���k�:�	k�L���d���&@���7���#����i�J�fB�ƶ���'�.?���uV�t���a��j��XOT:��^�zoe @�Ϳ+�v�m&Q�x잾4��>۸lL0�XE�C2:%p�Z��6��['B��V�}���*�7u�^ʄ��k���*[���z�=�Rq*���a��i�e�ވމ� BUv��>�d�-�;��G�x��+�i�'B�4b���i[R��?�����T��I�x)lHU��'��86.��,-�\挬��x�Cl��Ȝ3�=C�T۽~�k�aj5A;?�`U����鵖���\G�!����u�U,T�p�9�H���;�0������H�xy(늑�2û\\��|���k��z�Ĝ� ~<�syx�����[ꐊm��~��G!h�	�١�-���z/VC��2�V��CNXH�'�Q���Û9�A��Qn
��MlȜṰ�8��.)w/�b ����7Jgm5�N`/�y��p�'*rH��1��2a��ig��ՁAQHݪA�f��stz*E�"��k2�L�@,&
��q�2�����a�)u�1�*+��^xs�ΣfϿݤ��+-[�1������������0/��H�s���z@\	�m�o���k������]��v��H�3��֊�B�B�+�_ �P�i��
P	,�	+�&��S_ϣ�e��N�����u'�
˱멕C���a�9;L�+MYb͌SX.�BQ�:�K����q�&��6�}��ýB��|a��}��V;2M�{(�D�0��'�[�8�4�s����������3H��Z�!��VPiV�5Zf9`7+��xY�-�W6�t�+�|B)c�[��J�p{b4���q�,x�'�F�Y��x���覔@=YN��{jlTF|9�������(<_��m��-���Gzٽzs)ϱ	��.��� ������;D	@?��|�b\yS<t�O$֚X8�yK�F 
�Nj6�/���E�vP����唯�	�<e��i?�9���b�M�pܗ�b���{f���'H:��$�?_�{d��ʲ�T����O���ރ�H�rl�֜y9��1��X����}B���{eG�I�:c��'���v���tBv�!O���ާ�=d�|9��{E4q���{�E&��/�UQ�)��m�#��Xk�N�v��?��(,�� �2^uy� ���`�)�y`Y��C�1��c�{����|�p޽<��+�]��w�"�ډ`pN��j"�罳R�{�=�*������ ������h��a:�k��[��wk��~<=	�����ȝp��,�rfK�gXgW�R`�G��|Ѐ_���ghˊ�A�*Q<s��V)V��!����Ҭ﮹�.��~5u�}WP�5WB8��iWI�`j� ���}Қ&
r˘T��4���uI�
'��>�~�µ�Ԏ)߲��~�>U^aY� ࣻ�Q7��N9E(X,�B
Йh�U�A�[��jcoj벐U�m�0U&�m�ST��1r�y���w��'>���՚�0�o������_k�}�-o4>�H��U��r�i�)�Vф��y�}P��
�[b�J̨�����}͗�O��>�Op��Bb�>�6��.��P��S���K\����R.��dI�B {�K%i�/$��=Yo�s��TP��L�KA+T=�n�P�?�:m�~��ur�6�J����X郘�n�������l&�U�������3�?4���`�ϵ����}�9��&�V�	~2�˹�,�F�J�X���:
Ǽ?ٟ 2�V�p�lV�ಕ��`�V���}��7bn����:�fhu��S�+2eA��(߀)�yNVR�#y��o�9���<����g{n�je��>�b�z� n�_K�B5����I�r�fMc���.���7:�TDG#d��/%t7bln�/�R|����x�"�M�ђU�\�'(y���4�+'  }>5�C����&�$������F��!�/	�TX[�;�U��C3���Zw�P�T��¥�� ���BK��Eج�"�����`/DQ0&Ӕ�LT����N�(	3E�0��Pd��2�_/�|��BJ�S���y�g�'��XbE�kj�+͵i3s4��������i��4�����:�VK�!sӏ*������s'����4���>f��1%f1�/J>�{�<L��:���:�'{���c� =�zz�k:ц�PPc͇���U�h�w=[���f�l�~! T�^.�È��M�T��T(�'�l�T:@e�-^�
v�	�"���i)���o&}wρULl��x翮G�r�9�7���.&����W�,���ݣ���������L�N�Qq�3c���葀���q�|��>wTK{u/Fb]2�)\{��m� ����t��^,���T�g������j/lzC������<��I�WD�YLt�9,�+4s��<�Fv�]6ԥ;&slsG6�+/�^���oͮ�sS�������%7��*��uI��x3,���{���łI�Mz27W>5�vqO�Ql�)7�d�-�(���;o�����t���P�X���w�����s�ù�3�U�			d�܊�H)�v��Hc� ��L�������.j�:�=�Bz��� xł��H�d
�2t��wrs��D}�x����
�~P�|��B��/��d爸I��."�{��tP���Nm���l��+��;[ӌ���P�Or?����.���
9Hfՠ=��'�4$�x<c���S}q|���e��ٍ�2�A0�E��fEc���OC���~ѳ�PG�m�3��M����]6�5>Iv�g�tM��� H�ܡ� /jɡ��쫻9	7��ȕ�Gm�j#���@�/���Ƨ�@r,����a���ɜ�	|�����16���3k��~oך�*S��Z�����m+�H��Fp|ƀ�c���6m�K0��K���2r�Xd���i�ǉ�5M�LH-�f3�j�w;ݩ�!���1�"R�2�?(�[�(W-E�w���U�EGB�e�NZ�-S�\��잆3�Y��0���^y��;iApj���6w�R28�܌&]A�y��5�>�d�z���g����,2�b�q0�-d�b=�j_�D+�:�����i��gfH�����$�7�x�m�Q��jH+*�b��:��@�A�YU� �cD�OU�D��u�[W3�3���^�(v gms�ްG���{��B�]�>;%N��p�v�¸���!c BC>
��G�LM�e7�>���{X�$ӄ�X�,��GQ��4qqc�D%��&��^�E�?)��u���#���o.G<̲yE�n8��]��p��m��_����$���J�Ү�#HS��a����$wx;kB$�7c��w��-����d��*������"< *ԟ	����Z���"��w�D����h���-g��6�('UzΞ��`BO�_�u�l�;��T�xe+�"0���:��Ϸ��G���9��ݢZ�^_�Ү\�P8�oH��]�3����_{}}�t�L�%Z��	V��d�h����j���ֿ���;��!�~2�Vo��#7�F�u(6�y��D��Oc�wo~p��<�Y�j��2���P#�����$��s÷��o��Շi;?#?

��@ԓzlp��^�k���)x|Ѓ,#C�s.�?tp������=�7l,y�^o�Tu���<mѕ,
���e�jd9��D%��h���(���fS�77jb�� 8�y�i2��2
��[X�.c�W�7;Ί��\}�����[|[�o��b"^�E�^׻{����G �4���*����ڢ@��frUvz�-��L�d������SX�d�-e�gͶv�{7,�x�,�i���bco"�\���3}_hR:��[�>�RmJ2�3�˗�8��:�Kh �b��Q��W�1��HT� ���z�4�K�E��N�C��� �W%(]��&3���Y��o}�7��!]R3%�(��j�"�o�h�Ā	����J�7#=���[�����vL�_�@}��i�ީ���p �䮶"낔�RJM��x\�pIV}5C�������2ޖ���	?pPl^d ��Xú���u�-����ko�R蔘t�5z�&�p]�DBN�mbp����cwv�w\��]��G�w��zK ik>��0S�p���Z�m���&a��u�g��D����N��$��7<�hf^�}�X���$$����%5�c��eW�3�I�p��zDt�G�U��QKKf_$$��ӌ�Hb�Ca�=M�
8_�\���&�d�L�Y�����j�2+1�ط�|ּ�[E�ߡ���G7��^"��8����U�����|Ps�qJ��8P�4���t*�b����U<t�f8Sɧ��~�	�e����~@�6Ϋ�@��Ë��<߬��JT�D-�x9�8��)�m)��p6�mrL�Yg�*�=Ʃj���rD(����UY�C%0?�>uh"P�6����a��9á��Ζ��V{U�G���c7�gA��6��/�*�$��x�B���6W�%)�
Ղ/��I�Ko�d��ß-�O)�Ex�Ea�-(���t�ww�� �(f̎��&�K������l���'����Z�K�3܊2�ڷ����4۾��1�0df��q��S���L��	�.jz��T�w��K#�+X#���k�K��ήĈ2��+U�����z�A����
�z2�Y��'���v_g�B��A{(���ۖ����(��9�ʅ�9[lf��<%�n����AM���ݜ}�zpH�Ґ.xL�
`�G&�t�At��YWv��M�8�!$r�7�f#.� ����f���8��{�D� �[�q��7в�̲�T��T��Ɲ����{�c�iv��B�!�M�����d�+fٸ��b����66�W�_/�R�ț欅R4��J#�mqK��q?������HS�����gI�+�
J@��!Z	?P���tw� 3�,'��>���"}Fn���^v�~ �n
��x*���l�ƛ�%���뛵x���Dw�p�Da1���-1�J��F���x�+�ZiD�)"�;Z��g�Ɣ��o"�O {�#�㺐u�A��\��ǩ�Ki\�R<"�ޖ�D��c�U:j�c'F>jKj#���ʹBk�/ޤ�׮�2���'���'Mw�?��玿r$[�!�.�`7o_Prϻ�֍�R�ahw�F+����;.��S������_s:�����]'n��#��`��k���Ъ��;�-��U��J�����b+��uhMZ�r�n���@�E~+C�J��ӓ����EU'�+�}�c�+A3���1ߒ��}'o�鑈KH���L��Д�182�9�ޞr\�`��\*_6�
�F�����d.��!��I��l�9����:�&��8aj��C�X�Љ�M����(	�i�O��������O�� ��J���L��4�S�}c�{B]��*7:6}G;�|_� ���S,(00�q2~1dd	b�̔���F#	
��H��^�\��^p�����&7`��[��TL�xue��r��X	b�,M�u���A�^iaݚ��2tU�c��=�I�bDB2㯸�ͷ����z��m���$�݂�2:���×���Ei����c��Kݾ��5�WG�ZMY������=�?Gmb�8��r��4+_9^#Dy�!B���BL�v7��&Ul�Y�pN�f��W�i�g��:&,5-
��ڢ�� Ɣ��%/2v� ��x�\��7��"{��7�Y�Æ���Ea�/���Q�K8@�*�J���lY���֞o�|�3��?����i#v���I�/� uܓv����F*�꘾���=D35)�"�5��P�p�~q��M���������`ZY��1߂><u��끨.�
��11�=�TÎk���C{ۛ
� z5?t))���|G1|�y!�i���` g����,23؇�q�C�E,��Y}�f(,$d�ؙ ���U�C0�'�U�~�p�^L
�W��ϭ+@�?����C����3��<�o��|����{檾)P��k��5Ma�u�j�S�x�X���Q"pw)X��	�l����]�&�آ���8��a�A�)hy!��`z���?���-jAq��_
��mfa[��\Uv����+�u��:XQ4a[�kGe��W5����\hƿe�,{�)�{��voXa�szF⤬�����շ�&K��flZ-�&����M�*��x=	fvbZ.�B�>z '���P�&�dp~T�Z�/P�KWD���CWm�fm~v�c����w��z�Wl��$1���u�~*�vk	���Z<R��NV�0����^��2��)�O�Y|���=ũ�Sg%R�<��aV��& ǀ���:�NǪWpzh����zIdo���I��{'ǽ�����<7���Yb��K�`f����b���e	n϶���U� ghܩ&=y�,�f�!��,J3�<�T�gj���ѥN�?�6T�.����Sp�5㲗�uD����&�hJ)	�b�x����8sF����__ē�� �B�6�R�+�}���uՉ��0u?B޽`H#���Ē���cΥ5D���69����1�!L@lo�����d<}Ϙ��6�f�A7�Bp{\����U��u豝���A� �N�^�۫X��Ȫgv`i�W��I{��P��3�k�E�zo3L\\J²*�K%�(�+��8Z�H4s���lsa�zpq��!�(��|�$T]C��=�N���Z�RZ�%o���4�l��\�N	��1�h3ZN\�P�����Y�Ԛ�ǴP�CJ���#i��i³j�`u�,����]x��n�� s����.���8���]P��٫3B����ms�A��ij5�9���:{�������	k���#��\$��ɥ�X�~���X`|B5��<M�/� '�t���?����Sw=�z�iD�?5w��+���"��i
|ܹ ש�on�Р��D�s�f^Ц�_�ѹ���3����^<��ji�b��ř�3�j<٭q[�
��یR3�Z��Bj�+[ݾ�����]#8��SC&_AL�:A�9��"W�4Y�d����m�%E �j��h֮�9�2Mq׆ڭ���R͈TW�S��B�2�`FX���!�3���(Q�����;wT�zW��E5�(ԙ��}Oe0��	��yUD��`*�(��g����+B�kEl:�Ԫ�yE���m䋐]�se�-ՏBc�O�t�{��]��ad�W��[1F���	���M7O�y-�{�QV�ϣ��"M(�H_�Al�K��ޣ���͹O:U �a	�ek���c!��_�aѮ�ȫ̈́��pϋ��A$�K(K�+�.�R��ż@.�m!�}�p�t�a\�;ִ��E��Z�������m��U�r��6ǒ؆D�a}j�A��Ks׊��q��֘�2��
�d���3rהN���j4A �E��x��.��1c
��9�F*�a�(���٭�&�H�]���s����?G0�N��	�7�nn��{�42���^�mi������խŕ�/�e�k�W#¯Vr�qk@�1.Yk�
.C�]0>뤒Z���3\*����p\*P���R�+;�	�����9Gv�BNU�m�e�-zQ�p/=�p���o�����評�Q��E�h��jVճ�ϓo��S�3�0T�~& ����$�y�P�::�Ѕ��j(��/F��]f�i度��h�ߙ�_����'A�eMb{��0�]���_����z���L�{��{��\�AN��6e����hꨊ���ڹ�L��S�U�<g�\�S` ���-��e�%}���@���6�D�mH�Rl�E�O�7��LUih9�U��x��
s�}#$����N֮p$�C��N���ha|���b��~?,���^�ؕ�͢�&��À��}l�g��s��=e�*�E��EԦEs�*���hO��(��P^�D��>JZN7���J����|�6�c7�ڃ��O� mf��f��Eˎr��͗Qk�Pc��/����cj]�4pM,���k�.�����3C��)ME��ͥ��FG�zj)]��=���<��/�1��T��Ҏ�؛���'���=�T!腡�5���ڝJL�n����"��&t�{LL�U{���p��{[ftz3ie�ѡ��ee�O�i:�g��L�"��[��FcȖ��mj�䠞��ŵ�TY�51�{��д��T���j&Ki#������e�
�x���\ֺ���$�х9c��W��h����ș�?BF��N���bk����	tBC��%�P��B4�h[��P8��l��]#�	�#}� p�%�[5ԝ%����P�B�뮲�i�Ss�Ge)��Y�R��{�`L:n�]����y�G�R�*�`�έ}����w[y��Xq�?�W��>�S>-O���$9��;�֚�t��>w(��{���P��]V.�&D�"5�o��� bt�|�l����V�<	 Ƈx�U ;��������=w��\��HϢ�iu�!��0��T����SI�WnTt��pnV�����7?[�{U�j�F1	�x$^�A/xA�>"֧o��r�Tcޙ:TM�/�Jqv��g;�8c�D����$D�������Gr�9:7�G(96C���f}�?���h7���x{��fmcH�נ�n$�g(�G�i)[�W�0��o���1.Jv�W�u0I(�X��{��}�������#�(�}����fyn�S�bo�}7���XQW[R�<�@�b������������s���,m��҅OA�raR���d��q�^f���3�����a��&�G�8���g�����AD.�^G������@D�xm
�Դ^�绌V:��bCE���1fl@�d���(����.R&i�
�� ��#�H_#]Il�7�$���|�},�pL6v:Ҷ�2��n�e�)��=b X�5�v��^an�p��b-�8#��Φ�N���ū<;�����_�([C��o��5㷳P�T���>�KKB�$���P_aY�w�b�i���D��$�M-�9���)w����\>v觫��K�@cƟt����~q��)���������{������qr'�;O�.�l���"c;+m	�O�X5
��kT�^�w�5(��A
�*�zP���r�8��jsw?~�#vt�QSY,<�&��w�^�_%�{����(�#�Z(��f�s����g�>`#�m".q�l(rA�/Ɇ�{�+ލ���	-�q��ֲ;F,'L�����=}���9��sυ���r`����F�|�&N�7�wAS(;:9��4�V�3�����V�~[+e\5��T�-v��g��K��}g�5�?,i%�7Ѹ(��Wa�&�P�"����r2�,�T����v@�rK��Ni����̯$�~������%[A�蜮����$9[[���&�hݮ�v�zi�:�b<�o��4�s!@����	or܊�F���F�N��E�C���t���y�ק~�:@���RBm*A�d�z3������gi��'��l<9�y;�g�k����Ms	��Yq$���D ��,z�\��F�ٯ����[�&��B=mYV��W�$�6'� �Sk�)B�y���E�+�1S��dy�W3��h�4 �ҷ���,�Y2�@E6�� C��n�1訏aG���?}"�e-�B�K&"�Ezo3����'���=D����0��b�	6p:����9o�K=�����fi �	����(��f�7�}D�rw��� ���pm� ��i��&:��� �tS@%|`�G��Ҫ��1�m4�H� D���χ�uS�=-AĿ��~:�:«��;��y�Y��p�V;�^�lf�� �����/2H��v���nc�F���a��KI�\p�`5U-ОJ��*튯g����mI�2<*V|����6�L>��0�?Շ挣��)(��8B4��L�Qd�9���9�5f*svJ�jw��>@�c�H(�.��%_~�v�^�ԽN\��߶����<�|5�?�"ޞ@@��ܒ�����B�ġ�(#���k�4�K����jǮ��D��[��^|��0��};�UF"v�j��$ڑ������*w�+2y����L�� i ��=Q^�k�Wm�0s�H�t��΅�yY�t�c�/BmR��xV� T)o�F>�uQ=7�L�^˄�d����t&�����m�µ��@nw޶����w�JvNz7<�������Ku3�F��
�yY}At��V��tg��WAܿ���[��5_�8θb�P�U��+c�6�U��Z������GcJu=1��Ϸdġ ���O���W�'�U������<��x8����Y��_��q�{�}�q�m���6���\��Z ��'h�M�gV���Īyl���2y5$]�C���h�$(+�7���?�m@�N�&�#D�6t}x�r`�$K/w�㸪Z�������e��A8���r.{Q�����O�-4���Ƿ'�O/ 6�5�Q��X�t��1m��
�PI-�@�8�N��0�+����/�sUje@�KM�}��Xhq|����P˨�������<tXr�;4��/�y��"�F�z� 1�+M�!r��jNr?���|���Y7-� �g�|9�����d�(����I�ԑic;���j���SiC��8��I]̽8+`��,�#�*T?6�rq���g2���(% ��{�(.&�Bj�K��7:�w��接u��$���ЛJd�p-x�M煦�x�o��I9Њ����u����������7�A�Ä�$�X"88	���<����5�� |�q&.O��h��z{�d�kH��d�퐺��'N5��%GG`a����q¦y?���`e�%q�o�e	e)�z�6@_/�D!��Yl<�P��Q��q��vG��œ� l,x�Z��� ���7�f8ݥ4S?g�-Ј���Z>�8�w��e���ܣw�i��ڵ~&s���T����o+����Qq��;/�D_�2��%�P���Z����ǖ��`D{s�.C�A�('c��|	�w�����φ���`� �-j�f�Ҵ��-�4B��V}��G~�,@G��b����0�o,�@�r�D����?����j�T)�-}��ex�-�ǯ7��C`�w������h
c%�,�5�8|lg�.@.R)��[�;�%6G��	]3���]ܟ����?!�����aU��j�?�3[&��G�â�4���� �� oZ���[��)�ݟ���\SL��p�9U�(��^Q�Ǻ�l�������H0+�1����i����:tU��q�iG���,��ˬS8��lN�p�ʆ�=󵭽�����q��c���x4?J2Z�D�{�q����Z�?�9D���Sj��NZ���d*��B�m[Bw�L4���G��O��v+�a=�(��kL�#��]�:�Ɨ1��g*��a�[���8��;^�ѽͼ �����ǹ;�zd�ޘ�@]4"���ix��'�o�&���D�i�n�t���/s+k ��Fɔ#a�/v�F����_�O�G�/������~srdތT��<$Z��8�&�2Wv�YnQ�/��x��n�C�V�� �D[����P�����A�"���1^d4�<&ܒ��}���Ï���U�q4�C��>&_=�66�0 �LҒ�t��UO��g��_bΉa]�)ߜm�.܉(Zk����/�v�Đ�V(/J��{��=�+?u�)�қrJ2 8��Aؑ�c�8�:�ug���,�HS�$Ds��g�[X�|�(���;h\�pb���/G����p��ţ���0���g	�4h��:	U��?6�M�6=.�t%j뇔̝�E�x�\ UK�TPa� @D���ۡ	g���d�ǔ����؝m��l�(��]����`vN�	&_��>uO^����x�	�`4 l��r�f��ʁx�gC��7h0`��>B�����������9��9�i0&��^ZB�i͙Gc�g���T@.|�'�i�d'A�P\e��s����4�=�G����{0&9�ip�4�|׃\է�<��H�˲��V�&^�!4�a��Rt�.���J��X9Ռ=�|���:���2�[:Q�#�F*3�-�!��Ֆ��	M�v|��	۝\t&�z ����v���?�Y��um.#�
O��K���r�~N ��cJ)������͘�4���P�6#z�$ڗC1fJ���7gg9��8/�3�̃����0��L��6�@�T��]��f�My�u>�&����BI��!{������ݰf��'�-�!��ƞ��8u9I�I��}��*�쬚o��!�ST흞��+$k69�MMF��n�"���@��v4g��{ox})�
K�5cesErs6��^��FzU����e��1U�'��W��f��[����^����v<\D�6n"Tx�6��W�g��U�(t9�)�+���-(K�Ϧ�H��`W��h9�b�oC��/І��G�[y|�&iJhBe�A���X��4�M{�mFOz��z��	4@���R�����Ok֢z��� �64 G�ޫ_۲&�my�fM]�7:����8sJ MvS�M�����|�MO�"�ZQ{��7������ � �pI3�tj�3���_�y������J[�.i�;D����*�~{�.Q�x��-=����� c�<�GL=��r�Gt'�8u'{��� �{(�K(��q�`����HV<��z5o�T�A���)��t䧻�mU����o�SQP�
���p�!�X�ߣs\���>(�G�f�
�i,��WГj�=�^�Ū�6^��Kxn	�Jgg�#3L����J��mޕ}�D\�r�D[[�K~��]��5-�D%���oXqI[�I�LMD�4ܕ�u%��(��(�Dӝ	]VC��!�r��7��z9W��j[ݔ� �H���5j���F�D���(�@d[f��b�Z�:�NQ�� ;P�*�=Jy�n ~o�V=���șO�X�߿2u
�E�~_���b�'�v�ׄp�rDE;H�w��?Kցҥ�(�j�M�r4pɚ N�E�0Fu`�x)1CȂW�^Eūp�ַ;b����b�R�'_�᱿R\�ks�%]gh5��%?�Cb�g5q,I�fa�E(��Z�,9qd>�0�G�	�sz��O�`��++j<d�Fw�jjǩ�0��vWTa���D�=����O�}-��o'�{(k�<6���sg�ڇjW���\����0�c�(�<��k���x�lP�c�^JO�70���T�/�\ԴJ����S��ЂD�@���gS6)
���a����KoDSɓ�1T�m�a&�#��ES�{<O�~*��g���l�����_ ��mt�����Z�hҖ9��b���Fr�r�AZ9��ؠ
��bͿ��Q�<(ˬy�rC�ɛV}MaLv/�dk�[t]�� G/��w���/�I	�l,�h)f�S^C���c���K�g���7��@Z��&\��?g��n��W�s��x}T7�P�]�:�avh�[�,�\z�^�e�:5P�m�T�|��z�I�*h�����FV����� .�M��M�7G&:��Zm��i�ś�ڶ &-�$�Ι�� ?����|��dk���7����PEJ��;8Ă,����^w&�wU����L (�R����Arh� �P��N�kT��5�a7�U]߳���I��.�	���
ӻTn7[?#p��Ӌ���L�]�ˮ�B��G\CJ[6���T��U7�ܖX�ޭ:����
���T�E�X�x�v,�x�	��uS���uņ�c�	��-���t�\��v�ы��=Be�e����g�h ����E��8�$@�S�|(ܱ�EE��?k���gP���Ű��ǆb�p/'�و@?�BZ�q�5����
[KO�~��l����g�I�j���R���#��ѝy.�$b��t�|����x0ܻ��{�Y�� "�B���iM���A�Z���;T;����(��;��48��g5��\����MQ��͑��1��R7��e�ܴy�f��A���&�E��t��^6��4�B��͌�!�+]t�;"��"�:=��9 ��N�;�7\+v�1 ��$���zYb<�Y8�aI� z��0�G�ۄ�yDH�;س+fo]]A��)�/Lb���v��D �����t�@߲�H�[v�~�����j�����y��÷��B�� �_���9	Z�麛�(p2�_���?��d����q;X9��eBJ�lͣogX����_��%O��N|���SJ�)%�9q$�V1�u �C+��O�����bl0U���~�ZΛ��t]h�����b�v�`K v�/�	�EFX��g]�~r�0��*.��CF}��[���:`P��,���'a�����H�����&�h�cc%b�<�������-|S��������W8�Z݄�`X%.!9�#ҀMo�,��ɇZ�Ԯ�d��wBE3<���يBjh9�ɦ�_?����\����R�񙼹L�=b���`eڅ��S`�ߙ�6��"č�bz8G�w��)�C��o���_��%P����n˭�� v�	�u�ʧ��׾,B�ϛ˴U��2.#���)�,�s�7��Pu�􉟪���H������q0Zg��.����6h��`����̝��3�U���&or�G#$��lfZ��o�p|~7�Y=�����!N��>o�`�nQ�`ʉ2�������R��v#��U^��!ps�[9x����y�-{%��
ߘ@&�A�u}�w\;p#{�ג	��d]�ΐCI.�~��G��/4�&�^�^��:���R��P�c_���RFmy"c��:A�����,V�~N��&�:�L^�ˤ�$�C#�T*�`�\>(��c��W���I�57o�R��V��r9mL���%��F]�� � ��_D�N�L�q�>_�Y��U?=Du��:�u��*��!�|3ܔF�1���d��w�U�I4ͫ���Ec�EU� 5�<T��Dץ�?ŖD��n�wȟ�nr�Ž����a!��� ��o���K���.��K:AF��;��[��9����6�`	�:�~��D��?r�%��c��(
ii{,���H����`I�.�ۀ�f�S)���8d'��sï��ɱ ��͝:
�W�+Z��(AʢF���߱�ˆ��'�X��b�*��4��J�4 C�E�Ľt:|���£}J�H뚦4
O	�p��n���V~�>�.�6f@
����=�P�-SK�E��C��l�k$��N�t���5ep���AC�Ƽ�\ug� �~�L���xG���'���H"�&x��t�ך("������	nޣMd,Nj�}{:iMw�N��CUs	'.p�v1g�@���k!�	/nV�|���NE�c����'�)p�o�Hv �j(�V>��z�%zV�O��RN�:{3p&�j6���E��$����zɱ �GGi�`�"@�t����J��� �$нC!�n��ڿIaȨ�K�n��� ��+��R>�̵�K��/C�ׁa<�S�`��0��ggO�Gz��NA��]TMk_9�:;�6-T�+�	�Hj	kuqJ>��$Eюae�������8��j�f��N@���k���
�h�2=���~O�d:���q�S��@�=aG�u���L?���y,ݵ���	��4QZj�Nf��q�[*�c�!3����fPv�}[��r���`�(�Tɰ�8M<�ao��e�����է�ZbA�~W}40^:�hx�Ik���QeZ��n��^��D1�N��ӕQ0=���ʹ�4���_����sP0l 0����C��~��G��+h]�4�B8�$5�L5���Գ���"�<�~m3k#���pU������\�K���zO�����mS3�n�9���53=p4Y3H��#$]G!ԑv�(�H7x�,i�"�����{�~Ym�"��� �P:g��(�Š�����Y,餥N���]�pD����zԏ�q�v�	90딞�{"n+#b^F�E��z+#m�4kd�X{7j3��
�e��?m.���+%�9�[��>!5���QL���U��u?T����N&x��X����dB��'��[W8o��f��{PI}�(���~1D:�N���W@@~h�������ǔ�pT�+!xq���\����Pl���mM@I�Z��7��N�f�o�r��aX��;�ʹ�1�1N�i"�A#��b0�{5���~�+��Dٍ�ܶ�F��*���i���� 9�d �f�ܬ�<O�P9V�@��_ʈ��/T�<
;uU��?�{�9ۺp��l������K������/�%�.z��a{��q����s��&��43&1�O�Ey 5!����W�ę�(&OU���*k�=��W�DXI%�Lb+�i�۠�q��e�ΊKԗj�#A����
t�Nb�M'N��Ver`kw�Zl�㱙���e�?]j�as�i�r��J�x����D�@�mi�'�lR���x�w��g��鳏2�D�rm�j��C�7s��c!E�R{2�!���Ń$���h�0FA�L!6��;�f�,ǃ�ʼ�RU�� ��s#�a�?�����21^Kf0���I�x�w�3�Ȗ�`���Λ���K��ѱ@�9HBQ����`a@��٭U�},�UqV�,Q�x�t�&���9@�?W���X�(:I�'�J$x;=�g$�U����H���E"�͛ae��1ۀ��"o�$�5N�RP��3V��6>{��I؆>���>ÕM[X�<v�L� 9Y9)+�ڕ���?!��F �"t��Qi!�$믂o� ��2�A�l](��Я�(�
6�G��\�q��WJH�)��">ͯ��:G����!���@����FeVE FSh0C�j� �Z��o��wvTX��m�-+�w2�u�33�s`��r�n|�͋��5J�pa}�s
�׉�ם������a��2��%�͒O��-�NK ��M�� z�yJDv�c�D�6�븙#j���������9��Ýӫ.�[���"���d�eȢo;܍��W�Սc!�g�d����bX�jfԺ����|:�����QJ��Я� ReDsٰ_s���ޣ����(%��,	�<R����W�[¢/q�k���ئa1���j=x������ -1X��{.�k��^�g��L����6&}�����C�+9�{:�5ƭ��{�,��yl��*[�|� �H��g�S�9��Q	9�Wc���ْ��vh���%��]8S� c���/h���|67�Dǎ"NPf~�]�D�$�F�7�j]�8oY��|��>��,�l ��K7���{��Qr�xZ� �������ѳ�E��v��%5X��7}�_K/<I='��i`A��8ʠ�Z���7o�;�BRA�m�"U2��Q�[�z�z~=��Y�
�f�GSOLZIC������%�\��^����5��+o���5�]r�DŠj{���υ��xD>��+����B���(�naK��7dd�U�0�q������v��f��!Wd��s�;�]z��"8cR�w���(I�k��`7a�ִ�bѣ��L�~rd�r���`�vk5����4ng#���]�S�u�7����+�`�Hj�'n��k$�uƜ�>BV��{nK�ϛJ���d�&� �p'��l�Q漆�w[�EjJ��<��׷���-�͊�?U�n�;,��{���aB
��kȼ�N��Ѣ�Oiwvwcy�R�ŋ&�1j�@I�$��eeg�;
amVaD2��&Q P�>�V����Js��&!��7g���,���e�޶���'�}���D*�e��k]�����7h�^�,�,=��^vKƹ�j4!��s�x�]�MC�k��,u|�ںw�/���Nс՝`O��8�B3�]��iT�~R���;iY�9X(9o=�h���M�j`�=ň��8��B��T���1��U�>��=#�#t����ٺv�Sr��t*�����6�[����IA�>�PnU��RLb��ba�H�C��#���f�|��~6�����j	��6%W�>D�ٟvFϱ��K[�z�����p߇�ی	�i�$��Jd��W��j)���J�4p����ɖ[$g��_�ڑsV �����	,8=@o	=8
3�F�	ô�ފ��<��|Pk9��U��+�5�k�B�Vwa'�>�̳T�?x?��������_p����*�a�.b�P+_ [\Ȃ-AZ]y�<�m4tD���(�Z���}m�hMĀ�!�z��| ���R@+��r��|���^wTr�`
��c-��<4�����gqƩ��w\�������	��/����2�����tor�+���۠�([��t�<�j7O�9�U{L��y?qn�2�����%S��3VԠ�<���v��)p�(��=�P'�$4[^�-�y���Y���i�	���u�>�A$2�ݔf�1��&�'�"6��UY,�.}���L��Skr���9hԗ���c�_3~Hμ�]� �F��B�,���ޒ��|PM6��vE�D��Y,d7Vٔ����[L����kND�5��n�BD�#<R�����H�T�l3���,��.d�w[i�!Kf]\��U8����n��\��=��6�T�q�ֹɄR��ت�J���Ҹ}�,����s'^���KP�˚㗆i�ߌ�Pᜊ.�u,eq��K4��On�������ت�?�a����hXO��S5����W��C�&3J��ߕ+��� c��x,�ټ);S�oc��1Ǵ�+"���x��)���B��"lo����t�"�M��OL7��x �٠�d<p(g�ȂP�}�T�.�/`�T�k���ǘ5���ڼccLJ5i�|�j����&V��@�(F���i��q51��at�T�b��Q��`�sy��~�ɉ���k��&�j�ˢ�AБw���"׭�ɍb�ط�f"b]�R���0M9�O��������
��HR3M]�}����L+�z�0S��=\��q}$fe,�t�,ݴc��(�{�T�������4@�W�6x�R7�5�!����i�OҊ�.�%pAܧ�8ȤxiIC�}��w%�B�'���T�T�2�F�a�j H������6�>�E%�2������^̙�"�ߔa8S y�m��7��{�+��`@H��\�#�[���~���{�t.���n����cļ\J��,����FU)@h�{��ҰCGH��41Y��`��|{pVpȭ�}�<�¯�pbI���G�t�	��Hy���pefY��]g�,q��BlB��v���<��{cfD�cmM<FR�Ɵ���J�
a����Ů��6��Y��e�	��{:K�>�qJ��,d�'F����{?4+q܉�ً��H.P�P�����K��NЎ.`t?l���]٥�%|�3;��1���<�1�;�M�X6��ٷn�=�R9�߳C¦E��Ո�Ni��)
���C!����C�I`�2�m}�3�9dDdlC}l���1�:`#�R@ j������|��u���F�>��4B��X1���BD��Ά��8�bU�Y1U����%_�BX�*��s����R3čo�-}��4�?:7�����d��SL]�ug��0D{J��¼,Zt�2��X���o(��Cg)dLK{��F��}v�|��m0Px�0� -; ��&y]�0tV��������DS,���w���:�$ݗ�ddK������;���r^���-7�lN��L0�}u�U\b,�	�G�>K{�֪�_{YH�)�ZʼuU�)*�bԼl4�t�����B\>������\J�wD���T��Ʌo��M�p:D����:Ak�vz�L�5Ĥ뼬~z�3��8�t_.?buld�K���j-�#Z���Iڸ�h��%/p����G����b��2�3��:.��f��ʗ��|�[�(���}=$pPKQ���~�B��	UX8ޤ�kHC�=�W}jdO�y\G��.�x�*8��epl{+�׷Z�i�p���T�Asc��ĚV�NKO�& }.���QkV��R�W�L���u���܈TPZ-�XuL]�{ɚ9՝}����C���u�^�
nADNB�U�B�=�mM���e��i��=7�|-+?Qy��M�0v)����l��`�|���Wނi�N1D��=3'�C�W�%�S�U�<CqW#��^|�F��/R�D����!�R� z5�B]b||�DXH~�Mt+���gݏ;�����G�ߛ����1L��R���A���hN���C=�"|���"DC�m��#�Rj�yՊ5�����gN��<����>X�b=�j�4�'��}�D�N~.9���جqܲEM��BL���L�WN� �\y��u���)���\;��dQ�㢃-8Џ��Be��^m|�h�{����:��-fc�7��y�7}r�����̐ů�^*s���l�K�����>��E{�ݴ�J���j$6F�R�i��ІqV�t��;WC���΂ZH&�h_v;�B�(����6�Kˏ�*���}�t���%���C�Y8X�ByZ=�?Y�ԍ(��L.���V㗃���e!��{J_��F,��=����"�"͙���Fw�@?^/`\l$d&�H�s?5E�� �N='��k��<��x�% Ԭp{"`�M�y�}��p�h$ �le.ŉ+I]�fLW��M�"�J�M�h��d�[��(ZkU<�}M�|0�}Q_O(�����J�n.I$T�t;�ue������Dm����D%M����ș���y`5�ƭ�V����!�&*iBg&J4�M�6�W�\=>I;]�+z�pe!�D7Ǔ��45o+��v�P^�E��GF4�Btt�*�&pB��B'Gt�IL�%��C���B�
�i8mI�b�t=��j�hp|���AtŁ=�
ۛDK��v��$w�H�k@�:���wt|<{�l�_�Q�WӈQ�"b��nW���&���k��N��RL���Y�.{�A���u`3���f��Hz����b ��S�
��r�w>�|28��P ��a+��w�����4�XJ�oZ<>�]m��ux?��� ��h�/�_���:���ߠ�k~�����δ�/�.H`��*��=/����Zo�ְC�S�:��K�y庮Z��1q�� ��ʥ�4T7ۯ����	a}p�9akj"ͰM����E P&�m����cK�Os�$�8�}yV�<U7I�HV���������r�K�D9Qm1���T	��O��}wȥ��:o,���p�?y?��x� �?NT���[���f�{p^7���;q9WX7r�Y��U��h�����Wh�i"}At���~���5P�ٝ�,4$�[Ɋ6�7d ��=s���1�qNE�[�T��a���'�Ƥ�63��m�>�3;��W�R�%$��v��צn���mex��L���M�8�Q�cpjƠ1�-�X���C3���m�Z���V(�a��uL�
1��6���ޢxy>�@�c�~�3�~�Ҏ���/i��K^�����z:����[w�6=�O�]5)��ׇ��Mv@�l��Vf1|hw&�� �{�*k��SV�xG)~|�����2��r��r�+���_��TR*��x�2U'C�o��[hv5%*)������a(|Ek��0V�d�B�˖���Kƿ|DP`]i?�u e"��"F�ڪ���^�z|"�j�L����{�^PĿ�nq�3�$ؑ�އ�9:#�Uh9V� [ء����I	$�$sҎM�aN<OH�P���>Hn^c��y5K��I8��sF����U�A�{�n��֨��^�&&s��!���P8�?e!�^ΐ>���gD�-�ɩ��;۷�3�ui���{�Y]��>�yb@z�W�e�@9��B��Ew$Xnerf!���g�=�"�'t����Ŕ���M�pT�wߊ]��O#��Y�@:�{�8�qc�}7���+��j��{���Y��l+TjpkNo�V��L크�'G�-i��� �|��r$|$�yA�+78�o�3te�v�z��#-��=����@{[t�(p�H~��ƻ����5���UTC��<4(/>R���^�$�*;������rF��_��~����_���C�'���:��c��p��H��ƽ|� ��a=c�1�G�[(������YZ�M�[R����O��,[�
jr�2*�}r���;�{w��׶m>\O��P%ZT�ԫ�W�W�DD��bV�\���\�w�,�D�2��@Q��0avK�k���$�'O���1 +</�������Wq��@y��b�01	�b����dY���'�:W�4.�s��W�v�s�.͕���#�MB�O��=��֘�|�N?�����n׷�pJc�F����13�̾q��LdfDA�BPW̽����-*h�w$�L�ogγlG��{v!֊1\I��Y�����<Ў��L,~
�T��g/����A���°������l���t=�A� f�c�Q��9��U�eϬ��@�|�m��d������H�slI}zH\�n���ʭq�KRJ4x�����;'Z3���L =JBg�Ą��>Ew�٭���$F�s�S>u��%�X5�~]'6ƴI���!H%;H�uU�d��YU}����k�Y
���	^&��aW���b�IXmV�ęP�u��(f��E���z8{���J��Ļ�!����#����綉��T"q�5K���RA�!�ܗy� ŐFJ�3�1���.B֮�J�[�[�Sqh�^��{��]�ȵK���kO��n�n�0�>V�+�:�K�3%ȷPJ:IA�N�h���J�F�uwL�x�Y��\�#r�'�˲�cS�379��,U��2I"�?�yx��RI~w4��0=���0 �c��H2�`�dh��r���6�-z <�uw3�Ā�Ί���e>���%�qZR7,�LT������M�U�K*D+YR~�r� ����,m��c����eY�$�DZ�q�"� =��(7a�zP��9���h�x��o���E��eb��6D��b?���`���"3I =��Н�hLSQ���Bs��ڊ ��%/Ir�XR�4"�t��x}1�R�nv�K���x;r�}�*�V\߮����g�=�8�P�Z߄^ *��q�˔���w]
�	Օ�J�He��*(�|�M�f��r��yԽ�O0����GFK��ڀ�|,k����E����yT��N�у�awI�됹�/;=���D!>�fҸ��J�Q���ʈv�H~:��x��AQ��w	��6�sO7�j�)o}��(���a��<��|д{N3�㛬����x.�:EgU�f��S3�^{�2��[T�(:Iz�_�HzB��{�ݒ��͍�񆕝���BX�zM>�M���n�!���D_���{����-ws�X�t���D�0ϲ�C�-�"�Y98�(l�܌Z���I'�"�=7����;���c��	�-�Ի����T�t�/1���8>���o�t���lU��Ef��I�x{�^4�Wf��_�1j��@��R������=a\����|$0#��y�R�8~��Cy�Q��1
'�:('�bS����[�2QS���;�yHvqs�U��ۇx��2�7e���Z�Z�eA������L"|c��h2'�h���8����\��#���Z<Ņԏ͡�mZzi�`�>��0�ܗ���ұ�0oq2�S����ʴy�r��G���"�:����$(}2�m"�I�IE�)��M]�񥬤�e�Ϟ��&;�P��[ݎ�Y�Vz�>����[������8D��C�D�6(���:��yF55��)���};7���ⴞD ��zr5 ��]����9�pn�p��>4����u(ݴ;[,tdr�����U�]z�eA�~�%>�jM���P"C�z�>��t6w>��7�(���|8�7y1)�d]�m�"!В���{Ö���k���0"_�B����� �I�����:��p�
��ʹ �1%%�&�׈륲˨���?^�q���C���b���jQ�40Z񉕺��+�R���䏝sP0�v'��VSӭ��eEXjүA�2�>S`L�Z�B�@��1J �i���[yTH��h��Ym/T�T����$�IF`�m�X�}]������Z(@�jP�A��:�M	����(�q�f�\����j �e�೦�='h�X�������d�� �JLBg�Uߒ߹��K`̾��C�]�PbQH��V�o��/W�J!r��)��7��s��1A*6�����2[/
&6�혈n��P�k$��Ѱ��ml*���K�?��1_�	|�Ɋ��L�?�g�O�/�t,X'$�U��(���o��F~M5G�'�\r
$�۲�(�~g�Ҫ�^X�N3��-��d���9�\���ːՖ%�`L�S��!�h�QH�z�(M�!6�rٛ�����O9���Z=(�T4�T���S6�{�m6�a ��2u� 5��������⬴nP��$�)���WX�Z����r/�[=��@����E�T�zKL|ϳ�YdYB
��9�Xڼ�v<�V��@R����w����BjB�?��a�#��4{'�qM�����@�ɝ�N�	m�,�G�k$[<͕]7�5����h�w`q}e�A;t��fz�z�bQF4X�ϻ]ǥN�D6&�I�!�&m�Z��hR,���n��_���m�u�勁�LT�}b��w������P��W{�G���b1�����R���&\��r�l�һ�=�������9@,��v�j��
G���,#�*A�a�ŧ�΃�s����#���ݍ�����n�������~�e�����ΣE�%V4��@����V�����Hq�=X�sA�}o�j��6Vc������	2M�9�j�|Ye�x{qu3�I�V���CQ�uK�l^�`����y����$��t���ЁBX���ķ �&�=Id!��yK�����P��1z�ݨ�PMk�і�	�7���b]��®|���7۪�X��<��LW>7@n��� g!w"�>�ulK�f���̠��3��=������"�3͌��V��eik~Vh|O�����+�>a�����5�  �U*z#�@��D�᛭���>�۫�R���oq�L<�e|	m���jW�
0Ʌ��?�,���C�&V ���]�A�T%�K���h���-d;���*2PP$_��2��V�	e�VmJ�=<R�O8u�gh  ��L2���;���+�^�j+�'&)00�!Ӝ�pVU)���\���ؗ�N�2�ג����ȥ�"G�u]��,ޘ�t�O_�F�*U_M�L��m	̰lX��]<d��h�7���|7�Bs�P�7o{�t5��+���<�۝���."�/�	�8k�t���z#�y]�tH/*V2F���4+*���=_�r���8*��H3��r�P}�?w-��s��|~�gJH1}�
���,�!z1���m=�t��e26h�pg�7M�_��c,�l]��Q�c^����Eۊ�-4�6p��k�K�L�sY��d��`�Bs�K����uɸ�Դ gہ@�b��+��?����=#k KRX���}�,�ɏ�X> ����C��O�l��n6L�k#�8��.�����z���l)ɚW~Fj)
��E2"�	�<�EP=�����Ί��h�}�l��}�!oRہC���a`ws�,��<���pZR8E,�[<zm��o�RS΁�w,0�Nlభ<�x�N�OͫJ�U��P�v��W|��p���U
���F��X����݅��IZg��wջz:�G���%׺�+���_,c �f8�zK+E=����P�����wz��)��Z�T����j��"wa6\�B�	,�"�$�1ϣ�j�4[EN���l���$�������a��M��=!.�9Fkt_0�(SR7T"cL����S���`���?s��,��E���8�w��ܮ���ͧ��6.��tf��jc锑M*�c}R͏���S��H�x���y%���Q1�҅C�nm����K���`|U��|[d��!Aɺ/+�i+w��s:-O�~ۨ�:��v $�d��Y����S�pBF������S(��X�+�%��!�~�%��y/l_]��&/��K����~��!�f2a-i��b�vƃ��V6�M̀�a��&[�4Y迖Jo�W��j���E��vv��t��}+06���x6Lm
��*���F��AGŚ?����b��CI�z�(�M��GYf���T����ÿ���h�^yD�&3[bKߏ �`!�3��?̐�-X{����$!�4���O��&+��7�څ�3Ť^��0�y	�4�]D԰Sh��������1R@�1}���x�Y��#��h�$�Cܐ�F"ԅ�eʱp�tB)�GZ��匌��@��;@��S����У9݆ܬ�'��]p�׺׽�AޡW-�wr��X͡y�q��d�#=D���E6��{qZ��o��ȑ/�8��GJ���}k�v�~@�ގ�(ϖG���/h��+��;Ut�>w.���E�(�Ir�X���!��Z�!��#�v7�h#�R�U��tg^(H5�o,�G־ß��7�dW��B�OB�1E�eGC���.�1M_:8��s|LWx%�%�P�����n��nJ�@
Q1�ǰ�;R��$:�<�MH���Ĳ�n�����
�Z�ܮ#Q�i�]O�Ƴ
�Sy�HBQ����C���1�Ɂ��8��� ���:�
��'��m����(DRܿug$
~��'	�-V��\ֲ�<�u�hHc6�|�;���aP�p#큺�":�(��`���bh��V��O�d8��R���qc��.�J�Q^4�	���1�_4FmEG���/Hc�}�H��T
t�c�b���Q�?(�A1*��;���y�������˕�HN/Vٽ�dB�V���7?C�4xh��!�������U�el؟�t?9�հwOh���� �=M��t��(s򓹜u���Y��M;��X7,{��\�P6�;u�O-�#�Î�����*��yT\)�GXs�/&�˶�S2#XGP6}y��4}egDw��C��	�"���04�k�q�7�����m���@4�:�/(}��M��˻�Z�}��?���A� ��RH�H�3��=,cM�[h���w���m�E���"L1xI.j1�L�¯x��@���B���p�𦴾q`����@w��bt�m#˅�L�"/���W��4!���8A�?�s�vw���&��v����pF�ܧL��R�g��)�X1/I.��D�P�x!Ż����|ow����9}ZDQ�W�'�����<�g�Ő���:��6b�`N���~)u�!����f�li�JS����|���������e�ovM�m4���޻��ݣ�w.6���
�_"�	�L�b��>߀�@���d-1r	g�F���!�Zs��Y�vT�=�bP��zp �e��Ch�C�7���S�9K$�Y���cQL�m������C=:��'T���t,9+i�~Q#ϰr���d�	����1�N�\K��O��=���@�l�q4h����t_�ꃀ�0���b/}n�
���RV�x��.�����jn�U,. +}��ݐY�3�NOʹ�e���b��H\���#�j�0���_�݀-������c�S6A���ˠ��v���;���/�ja�����Du��$�xm��\m8����w��!��F��1(ƥ���!���y�0��yr.������(��6��l�e0M#��g�����/¯x���i��35ɂU5�|�`�9��Lո�Z�e��|��4`��0%�W��;L��1�N�����K�j$���Q:Dz%��jՌ��5�������Hs �	,�CA��0�0�Ps��ɬB[�'.Ǐ�/0����6�KueA۫Ѷ�Q���.S�Rf�.����:50�ɹ�L�G�����C�[��؍�cZ+1����oM(��%��bA{���]���#�mc"��^E��I���OZ�|��J,p��[x�P9������ ��ѐ^�/d��{%�6dx���|�ɞvu�IѢp>����0J��!5��-phN����P�h��2�]7/&К�F��e���?�F�> ��"�l#۪]A;�{y��z��Р<B��g��h#L�l��W!�������p$���uh�G��A��5��bp=Q�HC�ji��hߜ$���&�^�9�o[�*��y��78�����pM�`�>
�ZN(�	�)���io0�5�;VlRe���J��C�:�!�!b�1M�R�T�����_0�[te�X,��M)j���[���۱�w�c~�u�1�n;\=H��2�
��[�QRh���ss��JS������vO  �B�4GO�(p�>���w?rgd��O50��#���8�pp�y��9Ŋ�
�?Q8ʮ���][�Zz�z��N�,m1И��
}0evF֡4�[ɒ3x?�Π#�N�}�6uFF��/�*`�l���9�$�0]V�a�L��8:��O��{f�Ć$K�&j�0D���FqN���u��x�!�{�s>�g�r�8A��pa��,H���qCp���1��]�j��t��wl���*�3r7)%/%�|��g \�6R&Ü�F�w̓����0�W1��AJ+�uq�E���DP��r���D�L���� �;o0hy(��*~ꇵ��$E���`rw��+6;�~���u|���K���nZ��܈˱/ ������K�f��y�C�3�,>WO���Q�us��A���AM�[�=��(c���v���������z[??C+W��e$���~:+�s�K��8�7k�<���fD�{S�-=i�s%����$oW�1�(�6�7�n�έ=ZFl�Ԋv�fZ*:k��W�� G����+}�&Ơt=%�kzѷr-w�W���sS����\�sxΥ'"�(��Vݲup��bҋ�Fa�"	z8QK7��@;�����v�tW׬X&=}t ���&xy��V��̇����0p;gEa1��}�3���hR�a�/�ZW:��S#k9��qh\S5ɚ�X��y�y�����I1�}B���G�m����Vv���^��ZA�F�=��M3�u�a�D�=��F��l�N��N���>�^����� �7�gƫ���r?���o��)��޾:p�"��:[�T��/���������z�^�^�c�ӯW��Q�@\�����ۤ����<������������>���k�P<��ĸ�	���^����s]X���� ���D�Y ی��6I�-��.n�4��ն^�7Ģ�jN�r�EC6Cq�vL���,5b���d�mW��ܳ���A|$�t��\L�����L�귊�=�x�ݛ`$Cc�>�1M�O�z��]v��7�}�}cQ�@�U=�(0^z����N~L���r7]=�3�נ믉��8ѷ��Er7J	�&�2�/�<�q����Я��xv���"*) cޙ��x=9=Q�������B1���ZۍFPs�S�k(������cW�#D���o
���^��鷇����LPN���86�V�2N�D��Is����sL"�t�\�b�F��g8�~;�+��c2�ABa��9��S�i.`-4,�b�)b����<�f��	%����wo%n���_#Hoq(��X��Z����%���ƃ�Y��$��ﴉ��ϖ{�s����ޜ�Z�ǡ)������JQ����E֫��:�ɱ���&���OZ+��V �lPvѹ�>����TAF���N7�:���/|-����Y|�P�����^�;mƜ0N�fL_W�b������C�t	�2��P�zx�ȁ &L	�d��jn�x�ܴ@�WNG$7��R�`�,�I��n�ցa�l���}ĵY+]�݂���Il*RYmVXɫ��$�U_X�)B_�9j�P�,����4 ���ZE��M�ы�D��ȿ	�����_Yg������i�s���TIi��I�´F�gN�#i�t��Y�}\�j�DQ����T��2����M���D� LL��7ee�����o�c52����@%?%3m�}�U�4r�Ծ)�������K8Ŝ>�ѸRqB�.lz2T�	{���)?���/ �b�<�U0᥌��M<m錑$��H-g�i���H��m0�L_u�s����jʏ�� 5��;?@�q�izM�2�_GG|�Mw֚e�2�`m�UH��V�N9�s>pK��'B+��KlS�1őo��}p�0q�ku*��ݬ��M˒ϟ���Y��2z�5��=!$<kP����{�K���RNr��PV7=���w���8�ڡ̮@�u�,q�?;�e@�+3Ӄk.��'�GI��ڬl��,"��ГHW� zLh���=Vi�rFX��{f�mY߱:o�u�?)��E���V�LS��`VnI�����%dң�}���0M�S�]���MeDo���f�0}����~'~�3�vE�i��t�q'.�M�#kM�ǱW��;�n(�閁���"��%��`�o�I�R���D�	�W9�6�S��@�m���J�����+wPơ�s�v�9t=^���S@�G9���Wu��BnGt�׷�t��I���zt��G���Ҝ$�c�f+ؾ𠒍��g'�lz�w��22�����,���=>q���?�E?�����F��,����o�u������kS;?�o�7��h��w�<ɇǨ;~2�>�w�zمu���<)�D'���V떇Cab{���?�75v&J�Z�w ��	 �d���͔C�I��|����lŖ���2>Ϸ�&h�fL�C��3��ծ,���%��C��t�yL��O<��5�����7�4`� ����#���g�S���C���J��2�%�ʑ��(IF���A�fLP�;����tCP7D��K�В�;������ �����~-���B�y�cz�|�KM��8"]b��9�Z]�F���"Ò[I
}\�䖮��:�K�\�` �\$$L�����]x9���T�|��u�e������:¶���{�h\ɿW�0�6 �w�D.%S�)v+��|��a�����xT��3P�}��Sq�1��3a4uu�|6���h�c�GZr4�Lj1�f_Fϼ� ����gL����jGk`�������y���v9��}�5>�l�!/dB`p��Ȳ���5�J�@5�g`�=rq��g���Y��E��Ph�@����H1������],ښ�$؜�����[i���Oe	��c;芿^�ݢ�d�'}��l��T�Va�]��,��w�|�'��^;u�"6(���ub��b4�,S�n=������W�|����[�)�+�͵��zP]���l�z��7x�*��-�p}�=�YrDku�v����v��]VHZ9�c��,�3���z��±�0o	W4�]9���")�S�7N� 莞Qp�M@s!�S�H�1��W&�6o���#|n�`%� �ϡ4Ї�ɭ��B�S&�]��w�)T��{�<�<ޡظ$�-a�h�G�Mc��y��S�U`Z�����sp�Zy<8q3bXQ_��p���@�bJ�߄��"��l�
���Y.�+g���#`6�DTh�^#�M�:+�5�]�-�Mw��a�F��^�S�� �"\���|D_�|����6l�t�{}�oF$t�n�`/(mm�̈́7ƭ�7� �ڱ�dct��B�Vuu��Ͽ�ܯ��&U�?mC��e����L,�2s������X��"�'?܀c;��IC3l���\�s�
�-k7m��kK��HU��<����g!f�0x�D�='_�vv��^>��%ћ���_N�����z�,;}�OR��}$Iډ������YK�-�uXH���t�ؿ���?U���D,����E������of#�6�a�_���y
�V���0�0�0�_	�����\3�@V8q����3�Z�(��i�w���#+���T�**���y��!����m���Gã��s��������Œ��*�!yAK��R��Uة�����BW=�a|S7a;�����^�8b��~���r\wI��?�\�<�M
�T���ꦐ0VU�S�R���Z��X�<��/�)?H]Fj��H��;���=�Q�ވ�,���&�
UYꄠp���,������.;wЋ2�&T�7 y��%�������_4A�c���O4�f���p��@�r��U�T��0%Q���;���՗��n���'p����q�`�7Ǎ�T���f/�["�]Z�p\�����jH�]�K��L��ͳȠr(�-�% 	��N_�e0�4�m���F9�BK92�õ�P�(�0��;�KQ%���iM��߳`I�|Vn��S��Qf6$G�F��������1���*SK#��G���N�-����3;�S5��p�}�!3L��6A����
�9�tŶ��B�ED��q������ay,�w�P�W�t��U�,��#�� �%�2��pS��XELW��)[�>N�3�BF	{D��:��&�-ieQT�J&M3������gj������Ї�2r���	IZ�cS8ەR��s�� �����<۩{���% ��U�6��w���/��xH�Ɯ����r�z5� �&:�"̒���|NHNf��B��M $�
�*���v����r�����@���x��T@�ؽ��p$��ACn9m�^�|��r��Z<4U�����&��6�vGPسa{T�ny�;��n����ʕ�+c�?yq�a���g�$g7G�A��5�2�i��`62���%��@�[3{~L)��ڕ��/�lG���i��!b�٩Rh2�]���HNi�B��D��$�x$쌃�u%_�X���yx�-F޳Dt$1����#��ûz�"�r�#�O�5�����4���n�*8.2�4����Y�_j�E�cf��^�f"yu�K6��k��e�euJ�+�{0���-|����T�T�~��������<w�R`���n�V�z�7�Ҫ�����*��5U �isDE&��C�7����	�¸I�ðA!��Q%�5�!\c�0wf2�/�&V;i
�P��\�J��.Y�uXJU��c�R��Ҍ���8e 6s�I7�q�����4�X��/zk0�o�1�
<N�ҵ$����Gd��>f�,[�5�G�7Ӑ2�] �ܷ�d��U����q� ^jPx|k��A��7�":G�Ι�'Q�:3�HA����݁ya��.�����k!���%��U���к��Z:�4���r��V}��%sH�<��+���`�����<�V�R��)�@x�(������C�Gi.IY6�%�֌�>�Y\�7=�\�0��n�����e�i_ �3��)(>m�[�	�լ�e~w�t�煪�.z�ō�;w�C4=�اGl{G�,$Gְܬ��*k�\�����V������mL	�I���r�z�����B���r��%���w�Z���Qs=�������<?�ǆ(!��'��ot��:Nz���o��?>i� �X`o{N�JP9~澧L5��lJ+8+w� ����U0�$i��W��%*ֺΞZ1�-N�F?n�E{���4D4�r�k�Ê�qb���T�3�N�6j!]��<�H�ϊ�_�-2��p��xX����N�fL��f�q%�ļ~���u����t������e�Z/۩r�vn���>�0�o5|nY&m-���=�Q�W�A���i�)��/�1�X�i�a��a^�?AE&#�QIv�)x��2�p���d������H"kC�5��ۍ��%�p�|=̟Vw�R̼9����,-v8!8:�ʣK��T��� �>g�p�'*,� K�B�@r�6��w mx�h�c7�*��ԬЇ���^���M$�l�!�/�@��[��D�.�3��VVǼ�K�{�#��5�����8c��HR�J��?�
�A�����X��)�Ǽ�{N�A�%h���PسY�F&o[�K@�ŵ�dۣ��A�N$j�yeŷG0>^l-kP��3�H/�?LJ�m�ӗ�3��E�OP�,#F9yD8 ��Q� o q�]�1��2P�Yq�C���:L�2�\�[
�;�%��6X�]��Q��"' ��3��C\(�1��siܮ]�uN�m�����J�u] ��{[�˿�����5L��t�����Hb*/�>�n�5�a�?%�3!=�:�.�(PM��U�maj�I�����.�,1Q�����?+_�o�c%Г�]Q�V��?:�UJN~�<��g���Z�KB8�����h���
�$ 4"��|�-���ss�i�Q��,�$�D�7T���/��g��lv�*�ve-:�f-��o�p��!�zt���o�A�c�:_�g�$;��'g <�nJ��dO�TD.Sbi_E�EiVj���ٟ`��3���QGG/�4`�I�%_u��jU����QmE�,b|f��/1���tM;��3R@�5*3�T�0���v���Gm�gȑ����AB�"\E��]_DXz�"?R�I�3vuz6~>��5Cߝ�[I��. 4�KW�Oy6s)L� �0R��H�63G��Y������#"8y���:b��{�#fK�"�u���fQ��~_JR��ENVeu��A���{0M�[���2�f���eO(��}-��h���+*�-(���c�{H`;v)�;�Z|�pz�1����ɳQ������f���!�ӪE#EN��P��V8�;|=�K}�/����_�+)�ɏ1$�fC����4�bQ`ڢI�x�&�ק����ձ��Vz1��{�����=x^�(�*! �"�6us�+���df����3
VT\&J`�2y x7�Ŝޜ���_��LyZ'���u��y2�qZH�-9�t}c�`�Às���2�
�1A��W���`�M��DXɑ�|7�h��	؋{w3Q��!*�Io�Ƽ��e�S�^_� �K�S�U�6�(":@СH����{�פ j��I�KD��V�s�	�Ɓʰ���c%�C2�8���eY����1�@�o�J��T~�W� ����9�0��-�ﶱl�ۡ ���k;��g�et����Ȓ/(��m�hE��
�&:��bj*���^H��"��:ŀ)2�]J)��]AK`�Nh�m������v	��v��D���ƚ��L�5��Տ=O�M��t�E�$%�O�R�hK)��R����=ةU(rd q)�7���#oy�>�Q
�#��T���ނG�j���qi<F�yڍ��G�}��lr!)8��e�U��`��V)H��Ԡ��FP���l;��op����=��.�]P��=����Hi�2�-�?Oa#;����4�v�W�� �����& G���w�6�Q�׼1�� u�H���B�P�-O��o�EJ�����*��m� �^Y��������z�8��ԍ}�Ʒ}�^']-{�l�BQ#OĎ��b@��o�n�$�x��j\���ي��rŝ� ބ�M@���܅v�h� �����7��b��9墯�!�5׮�y�̖��{	��6V%"p{'�KM]E�wj�vK�*��Q�}��ao��8�o�CJ�I��@f3|�� ���EH����o.RY}oms q$G��՘G*�ԋ���*�|tF�kC�^/�+����-�y;V	�eM�	�_���C���B�̗Z+b����PO=����ѻ�S��W��:q�[~����R�0ճ��Q�PE��|�[�ō�`��x�ɠmZ:��<M�@�a+���;��*��B�u��*���X(KG&�&�HB�`S#K�27��+ґ�]�ƪ� ���tun�<.5Є�eV�qK�'�X��q9��Dyy{MƵ�=�
�^�<�ӟ�[�ȅ�Gb�v�B���ou�oׯ�Hhwg��o����y�)t�H2��<="�v�_���b �ez9_;���X��xj�"-Y��Khm�$��j+Ԛ�y���H��a$��J�u�jq��G��û��"/uٰ���LE��k�%��(H��o9U��Ї����{:{����I��d�7��QuW��r���X�>���}�'\�^1��7��H�j>�jh�ٸ��b��4��DZ=���V
K�"6Z���� ��63���seeY�騵$�_�<���`L�|����)�o6�8'Te\��Q2׌ f�ƞf��7�D�ݠ��m�ϝ��T�nQ}5Ē�V�X�&�ɲ"2U�6_o��f���Sp�"X�|q[��v���AѤ���������e=���7���*�:>���4Ř1�j�f;�%?�㕈x]�R78�ߗ����K!��7X7]���&+����� p�:�q �g�1�v���i4 x6���R��ikX%L�_���W�g��X���Uf��K9S#	밅֪m�l�~Wc�u�q�E�<�y��'On&7�H�o�����=��$b��t���S~7�@�)��x󰾤���@M�.R7V0��0�W��^�\��(��؆4�ԅa����o�ĥu�G4�h�i��4�J4և/�nV���DH�#ś��	hYx�/-3���'w��apYS��%���ẕa�U��*xB̓�\.X���OXmg]�<����l���{nPh ����
t4=T�t>}�����B4��Q���-~��.������z�֘-[ �'�����Lg�Bey�73��dm?�lmM�z��J`� �N#0��ok���9���=a�@�hM8�Y�4��(^ٖ��&��ؖ�)E��:���rf!�B�/��}�s�wS���kYi�Լ�.j5�n�#Qe�f����;��f�W���w=P$�P�ln��@k�z�r����e2@�l)��	����g�{p�?�b��٧/!���+�x���G��%����P/l(�<y>�V�%J�`�[ZG������3<G`�;{S��ˇ��(!uM��_���M��je�	����m��Q���E�yY�D*#�p�?�{՝T��U��ўOũ5�|	6u����q�译�u�|���\C.�A�6�K��N�r�  !<LAID����������>d��a���骿�f�]���V2�aB+l�{=r�u߮���&@�k����a��S��c�R)��7
w�6։]K���	��v����=S��zۋ��&�h
��r�(1�+�J�WuZsx�H���ΡrD���RA,!rG���4���e,����������Hj�����)q�P�̿�ī8wD+���n�ΊB����nvD� 0��$�����K�!t��X��^�9�9a�������}���Y�GXE�HY�'.�����_�g�4iM�6�!\��5���@�U��ȱw�|�v�c��7�n��Jd K���D9��CH$��9����w����H4����~M�Qv�o�EmNj"��!/�ns2~��H0�R����&��C���k�]\����Ap|,�����Vɡ'_9�
 ᑨ]bx�J\���&F��%��n �wt\�tX�(C:��]ˍ�	0���0�-?�cwo�d�w%P�oOR��*ɤ����wߣ�1n'lg�!e|�y^�2�su��έ���Q;���%�? �͞�ڻ۹
v���Q��ή8X������H���]�A��G��'����7D-��M1�q�\jaH�| F�H�驕�IÄejDO�wp�',?���Yj��Ԑz�������c˴���9�T�6�Ee���$N4
q�zť>��#��k���~��E>[ao1]��=��c��YK�Z�ۣ$��(JBf��ݘ�n|���h+=�/��>�:��r
Np��&׬/��}9��:Ymr�=�}���~bmf1�v�ã�H�	K�a�,��gd��o�a�Ҏ3C�`[� N��En*�փ6Di�_���O���|��<�8����X�4[w�j�O��	�M�u-��ݕR���&��p(E�Ӄ�ڣ,ݫ_����BD�ߎ�( D)`GJ�h[�:^1��o��ll�?��]��R��S�4j������nk���p\`��izP��S���Ċ'�x�6�v������q����;R�ް�mSV�0|�uI�r��c��c�b3Wa3z(`;�"<m7T�56�mnI��#�D�ߥ�g�v�4�WN��4r{~��5�+j���%Kk�g���.ga�{���6E�P�0λ�3_En�bۗ���&���#�@UճpQے�x���[��T���7
�C��rLt�VI���s�����������		.!��zRE%�"�B3!������[/���Rk
rF�nm�Xg�.��#C�|`�\�
��"��s�Y���v�Y5�۹x/=�s��Bb72-���]H�J�>��֒Jc�w��I�w�n�"�K��H��Խ�N���[-T�-e��j�ݦ�I��_Zf瀣���J�>��5j�y�R [�;s:�
4�|"�$4?�&�dq��z �c�������l�Ʊc��#��.� ��-NJ� �s�cv�˖�z���%�XY�6U�'�θI�@��H�5?�	.X"h�R
�]%v	�b���/�Fg�Hݳ:&�/��d1�8��������m%C�����R�0�P�5C�C8���y��/S"�rdO^IVt�)�1�P�#C���r6�l?�}�I}�e`���tAr���7_�}���w����N~t1�і���������DVw��P�����	��1��vzG��>�X�n?�<ީ7��r����M��&Ez=�8Х}]T�y�k\2�-[ŕhҠY�
ˮg�-�W�"r�<�x��v����#T�%�5���Ow�������v51)|^>�zYR�~��3���bST2:+\���]D��ň4kɃx�%c�Pk��x4Xۜ(�w��y�*������i�t����)�V.�;��s����#�l7W߳g��#X�ʽ���ڟ`o����t�33Y�%w�LSF������p�� �ȍkT���_���|��H@?�;z#k5�z�J]Tp�\R�����)��2,LP��"�{�ԗ���_7�r���Y}�8�U��aQyƫ�΀�r����A}��%���p�E���s_ ���Y�� �o!�4����o�ܩ�0�
�$��"	�'o�0<�6:�N�/���{%@�J�<�ӭ���H�%g��נ�$�hq�jd��=tyes�Db���.e���m��\6? ��p�c()��.��������URIkeiW[g�uL4��P�կ[�Ž-�qI�Ki���6�~��[��~�.t]HnE	^e%��9�;W��t��i+�틍׼���D�q�>ptV��J>��|9������_e@S�Í<i� ���\�l��usBnD���=e LS,��=�Fi"u8�eC�$
�+���Ktş�U��#\���	Vx��o���C&�js%ѣ�������ׄ�@	�Š$�>�&n\����n������>84���؍F�0�?�?�eb����Np�bQ&5�H��ʪ�YR���,3����Q)On�g_ ��9X0�<��X���=7��Zaxk^7;�K��ܫ�Z�_�X�lOo���E�����.!^���:�4X���k93��v�S)����8�b�4+^�q���)sl��cɤ��38$��_� �T�D{J�޳p]���oO����\/�t��J��@$t�5��N���f����y��y��x�������P�$�@7��2�5��<eHF�и�1��\0��V6�L	�L��²�*u��������^)�|g�2!�}�!c�c�(:�v�V�)u�G�P��v7?�&���M$�H���z?[���E6.�݌�	H)]�	&����\[^δP~fM�����U�"�঱�2d�s��L:��?�^�tTW_�E0\�R��!4�g��w7�ݴ=�[W��T#�(��洿�,d� 0������� �{6�<�WꛎiB�ᇍ���yp9��%\�V�M6?�س�eW Zvdx�}��JW?Zg�z|�}t$
X;�|F����Z���ā�m�娿���@�������_���vA�L"y '������f��'ܼ~�@�[S�0�Vj2	,�#)����/]�	&�K�e�|'j��.�%�j��8�m�Tn�Ѫ�+a�p��x~
yE���7I����>=�i/�ꅠ�!�Nv;����j�>�'\�K�C��:���p�(�k��Lg�U�!`��������1�"�4)�L~�tW+ y��/�	AO٢n��!��(hfr�5k���
�>Ge~B7�H|(o��W��FD��@�[��.V��&��C����c�r���P�	ˌ��X&���p�Un�Tj�c[��S�����A���M��:D������e���r=};2�=@̪kJ��`Dj%+�'U}׸������Ҝ?oՄ��@`	�hk\��?D��ÍA�94��β��h����b
*=����W�/��xG��ė`7[�k��y���� W�x9\ϋ �T�����f�o5X�%�� �t�'���u�+XO��ퟣ$ ��j2�.�g��ډ���s���~ߏ���;��kZO����Q�*���!ƽU��4ͱ<�	lp��1�@�X�����c�񋡍)y��!�����X�GfO�oxgv<H�lja!5w@pԤ2\*���%��<�ŕ�)\�	�n~H$�s�r����6wDw��!�ap��ъd�7��d�ۮzz
Ѽ�i]�a��]�4���@;6��CĀ$�J"fH�Z������#sVݺp�KZBoe����1��i|��,��kt�4�����DJ�z���g)��S?�ǰ�Z�:k��-!�oȇ=�щ܏drM��в�S���D�n��ɽ�nsZ{ۇ��.Pڨ��d����Os�Fy8��q� /YQ5����(bx����#�n?�2�撜��q���0��25.(��ZR���\��I��5��w~pE�y���K�FO�u�'�n/�Y�ϫ�۟���Dm�ö��m�}��=^�2O�"��1+]B	BA|�.�ԎL��p��Y�+�n���	��!h[+e�VnBˁ(��ø|ssgA�-6���I֝�\Da��Kd����w���>��h� ���뢒d���r d�u>��!��y�"FG��je��X|� ��z�����ŧl]�Sb��Ñ������J'�������!H@�@i�\���z��m��Z�~Z�H�+'���×�%|� ��H»�Q�_��»��ls�Yo� ���g���2��������]��Ek����P�I�Ņ�cQO��w[���#w��������a^��1!O��y��OF��8�,
Z�� �m)�l`#���<B1g�@ l�]��?'�=wͣGU �����%�.� �6�+��\���}�2�FPa~b	�m�`�Bl��, P�4�V�V�}�����%��Q#���(- �%�~t��5�јOL9+�+q�%�-��,z`W����e�Tթ��p��u��`p��Q�>6e���//���-�J�t;"�Y@������Ge_Y(7);�d�'�1�&@O�5e|�LYѷ����߂�=���Wyؒ�/M��3�����
�l`�7�K�VD�s����;uS<���P�?��?��lw��mJ�NǸ)��[�!�FzT�|eC�xkN��h���9�$ֿ�"p�K��zTN�1�~q��L7�ո1Xc�6�v��ѭ�PG&��&���f�b+�(D6�nla�$��4���v|���"�}���5l�f޽|�Nn��n� R�~
n��Ƞ�ՙ�P�@\;��c������)��,�
f�G��n�����;uM�h�xa�F4-Ck���'J���A���|2OHu������G_�28{�]���"
G"����k�w_�����C�2�U�Nf؄��`<YȈ�M�)*���i%!��M��l�P!ei{�酖�ղ&��M�?���\���;�Y��ԓB3xo�Ww����kM�yg�a�'_3w��Ji�����B(��w���{2C]��^8��7�ycp����zr���U{/5U~��U������:��v�b^ҸH�O�7�#�$e9@���qgn�c���>����z4R�x�&�@E#k�45�kvqh��{c�]��<)�$��l[>u��+=�H���r%�,5x�Y������3�]Ƈ�?���gy�JP��rǱ��n�q7�ш�q�@���R�N�MZ�ђ1�a�iuH�J56�@4�0/W�Yc�>5���vWe������=�(x|���a�W�D�W��lW*䨿�	�M��D��c%/�{{7Q���U[��5��'��v����Ág
&��"�s�������$�{���)��k�2'̯���#�u?G9�]t�\K�mԓ-
�
��V��7�o���%�nCr��Ѝ�Y5�E�?�cN�b-Q�����S�_�aQ�5J��|����Ĵ�4�Zⷒ��F��Ni�e�v�o�#��ן2��Y%�����{�b�97���j����5Z{_�PD�c{��z�3�Sj�.�A�LQZU=:w��t�Z �O���z_j Ѐ�v�F;i�L�s�Y5�,:�p��ڪ�ҚA�fMV��M�?��qE���5A��rj��S�YxI��u���qz'O�A�?�K�=��@	�s̨l΅��p*��~�e�Q��~Sq�J�>��B����:Y�I 	�]�tkҘ��t�>ŔF2���Y�q}n����/�(��l���=ۺ���S���XXG&�)D�*?�˔~���Lf:.y�r�,� c��4v����B0+ѓ���i�2�o�BqɃV�Pχ��7R3�P����������q��Au�?[��b�K,������ �ݐu�e�|�Qm�(Ò2*����m�[�LHL����d~$Z��ڔ�[3�s�{J����l��An�����>��T��*�����W���u` �a��5��h�K�:�-�/��D�]yQ�Q��!�=lc����ӗ)�gn�6ҳ�dlP���`���$~��s��*���(��Y+MCSe�{�h������lcd
�b=���7��wrݷ�Yx۟+�v�e�@�hrv�&O�6W�gb�k�~��m�+�+?0н%^:���m��mg�C䬺����~v��t��:�v8(2��U�~��m�_U'b1�u����m��F���iN�n�0K��XH,�Ш�<�C��@h=wy?]%:/7�*��eu,��D˩~|�<R�W,��]^���$��!^F�G��q�T��.�{�	� #ޢ4(hg����mu/+��'�C��D�z�^@Jν3�/�:nl�$2��;5��� ��i�1(�*]|r��5�@�K9��*�m�A)�<�{���0rV[F�o��Y��
�Bf�R������ ��]Qÿw���'j�� �J� �fˋ��b����KˌT�;*Ԃ���z�Ʌ�_̠D���g�w�����/����9*'���N4��zLS��*�>=c�PB�M�vƭQ���m9[W���"i<�]7T!��)��8�X��j6ۡ�@��å,Xa�&�(p_�EX"V�d����*�Zѱ��v��QegX�9Y��d7WDf}=��B:0��+{��N�8p��*y�!;6�Z8�3�2;3s�K:�&�py/���iZ��D5kA�&�'lh�G��^)�\�%q6fٚ��31^��q`�kfǃor��o$�8H��P��ƹOzX��G}����)�v}�y�D�XǛ��FM�d�Ӡ1�.��CrWJu	o��j�4�$KB�D56���˲/A|r�E������S$S�(��b$�V�C`���-H��L�9lO�F.
Q'������؟a=�*0]Og��*r01��&����X�Z�{���{�j���^�@�8�)$�3_�����V'�1G<'���Hwҹ�����$j\*yQ�dq.0�&U�]��W9�tk	������H�85~&�?��\nDO�u���`5?g���wS�u�� x���N�&��)f�EW��%�`}�W�5=���aL���Ϯ����I�|��4��$��}.�S���#�)�%����	���F������[�@��hR���yǉ��3&�#x��]Y=*��UK�_sU�B���;߽�����
(�dpM�ޟ�Ԍ��)����;�c0��+]��2�S���䆌�}�-�O_��v��s�؃O�����޿z����}��u �
���G?��v�R���S�ymYL6i�"���ۺ��e*��A���hUj���G�;s�Q��[�߆�Ƨ7L��.:�g�|	�������Q���Џ��x?z�b%�[��gI���>uZ�a��k->t�iūqݥ�ilI��TT�	��4�[q���vΦ���BĢT�� ���5G�Ș6@i�Z�F���d��^���M�-6Ki/l96�[5�l�����=/�&Ϙ�=�C���"l���Z�w��ӟH��
[��u:C"�T�;:]��]'�
<5�F3�*������{�A���ɚP�V��#��XZR�D��B�k��Z"�{�J��e�9�*���M-_�u��s�F\Z�~LT_:�s:���F�Id�J�er	� ���!Tβ�����c|��b�1\��7�$L=B���,3��TݩOM��D�g�_\- �ݷ����$�]�?X���@N��w���op@��8�3�t��~�Ī�Q�|�����V�\�keS6c��YS�=^* #����A��k�y;
���
�`���DXp�#R�y�@��]����]_UO��pS  iRqgŭl����Y޺\�"�m0�n	���G�a�/R����b!I��d00�@Z�x{����^�-�슼��z`��1��p�W��}8����!�v�����!�����B���;��D�� ��+���Cz{扞'q�k���=u8A�3F�1�f��Io���+�qڜڀ\��@�����1W��=XB�g�۩d+0M���b�?20;>�`j�h��?�Q�X -��t�O[S��(q�[��y�=�����+_��sU��,K����!j��!\�ȣV�5��ezA������K��L[��g.f�=*�l�Pj����&��OᾘZ���w�t�Lq���P���$�*:�j�~c���[ �27%J	d���1��9W){g��wG@v�>��ܡ(uJ�F�2Ftfi�1w�v��EGST��Z��e/լo��Č���dg��|8�`�d��=�aZ̾l�����S���!ߦF�r0ĩb�d��:2�9�i|��=�`g.ڵl$�tW*q���œ�Tƍ�StpK�	vDq`��؀��96M��,�0�Q�\)T�~|��I|Tb<ד��X�Q��� �������^Y����H�v�hF��U���s�
8 X����J�@Ӧ����<�k�bN��3� �m]m�%|�C�q���((�0����4TVM������ӜC�rp4Zd���j-���f���$Wp�g�|4s��������^�0cyO:�|}ʝ۩C{��x��=$R���a�䇦�\k?�u]O�1���$�覧k-8
���������X�%`�H{+C���0/$�
�Q�^���ٻ���Y�{8l�+�s��r���B�m�	Աy��s^������zsl��ر��)O�֠�� �8`��/֦CP���Ɵ����#��$I�V4��>�+��]@X;e�y���AJD8��z��7mw�� ��2�N���љNK_�_>����A$�K��>�(���*Fg��7��|�p�u�%) ���D���	D�%w����!
�׿�x����a�p�L� �QM��y�h�bR@	'�HQU}?�E-�q�w})�ޖ�R�`�9��,J�Ț�x�����k�,�H��5�h��e�Sm:����Rٓ��� W
J�=��hj1}��8�j�F�Ez�sn��JZu��/
H9���@��2@!ep����qk��w��D+okG�z>qj](�kk���P��Up���!�]��(0�XG� &!s�����m���7���R�ȯ�u�ȬF1�;���x��@�QcYi�˭��A��)��2��D�L���,���`��^����g:�wpm��;��)E	�W6=\���BLD���`:�L{�r'�]�mKI�L��3j�v�n�F*!��z����惢#�X����-"f��b=zn�x\?ǒM�����
5y3�7T����0���3����<����>S!Ho�bK\��?��Fp����6^nӻ�KGO��ɻ���Wg���tv�o�&����F�Bӑ�8�2�|��;y_[��E:�t�2x��ӵI���q�zyZ4���5�Pw�(�toh݀ss����2�Z�؅>���ob3�vA��.P2�o��.ˁ���;��x�t�d4��?WL��>���۟���U̏���0Rr��v�f}�u�dWg��D���yu��L 7�m*d����"������5����:�d\����h�����.1�a�S{Uf��lw�e'w�J�*�^-H�A=M{_(�&!�q��<�ѓ}"mM<M�m�j�aE^O��hk�x�׫���=-岄.3[@�*���TS	R�?�B�sE�B��f�r��4>_���D�&�J�B�T��q�Z/��:��TF-f��ƭ��/���i��wܼM=35�*��h�i�M=1en9Ĵ	���a7�'Q7ӄL�{��7���ʓ�d����ʿ��xs�3a΄���1nͳ�&"��S�[�� ��V]xq`����8��l�A��9����]����
���y���8���s4�;�d��z�֟���y�����f�XIJ���9}(!��E��|�J�' (w�ֲ�b��΢'�LkBCȜ|̈�{�S��T3^���%x����(ȫ�?��0<�/��irGF��F�s��~�_D� �a�Y<��dҌw�%��g�����*��!��M&�8z�s@�ƴ�=��H����.[�ޝ���W�2v��$��њ�R�h�o��r�����%�3t����ŌT�n�vO�Ҳ����R5o&���*��
�)Ct��^,$e�����Fʘ��R6Ib�.!�ѩ	�`�������5e	���}�T�gv~�|s�oև]�ǈ�j�/ ���t<e���|�~x���Tb�}�(�I˧]C�M:]��L�Ɋ�\�՞���*]Z�� )$yY���+�J)�K6th�sk�Q#��@ǽ���o�}߅R��N)GG`�<��0Y�l��.�G���:����� ڡʧ����Z��(�P���¨��;�c��;?�m��5��g�h��mo^}���ʖ�1z*�����ce���Gje�l��c�7�A��a���>[��:�`ط`-A�<�ԅi���� )cF��/�\�834�p}��1W�-��@B�'��v��������5
d��hq��t(�*K�t���~e����b��1�pG4���}�����V��$�s��"} �½�{Y�~bY�e�6.=��5e}��B����b��<W����J��'V�I�@�i���6�eshm���(q���qq��kYBE�`�x�t����TO ��a,�-{!;k��b��@���|vՔi��_S�C{���v��<�����cZ�V���*���$ ����g�\����f�­
�����W˝�� ^L�����|>QXڹoo߽*/I�т�F�)��&�`P��쩩�el���j����\���@6�k�W�ڪS6P�����&}�S�z����*X��`A���h`$�ݣWX�t�|f�*�p���?�ln�B�{$��K�Z'����)L��=j���D�v��[M�֞%����p�H
�?���W��`R
���W�1��JA�gm��Q�{<�ɮ�X�	��#����q$�XF8E�O�����zJ���&����`�;/��1PA���H1� 5&�n}�g��y�S3��D�9FB��N�w�W�1�S�-T���ꃡ]������k��z��] |~��j���� ��Ko̻U��f��Q�k]AQ�M�|o�C�½��>�Ko�#�:�+��ݶ��S �e%�H�"��,���������?����e��c2��0� �Iƫ]S!��ޔ0."%s@�!�'�x��]�3&�3�w��r����I_�We�����8�@�w��=�H�o�$�A�3���d�&�x@&��7���h��{�OK��z=�1��@0vܝ�AE��C�ǹ��l4�9��n�l��<�_7t���\�6���F�ut�@�?� w�.,��i��dg�)����{RX���o��H��I��b�\�ٝ�"�����:��k��2�2R�^iBB��y�j�'��!v�{�l�<Pm<����,��q?�F:0��S���5�t��{[h�?em$rb,��<�Rȗ�U���=�j@W@�qzA� �	�,qF`�_߁�?�9�%i}��+�khp�m��YWR�xk����#t9�_�w@�u�N������$�`�� x�1���0���ۣ8G�@��>_��j�/;D�q���E���Ηq�t2�m{�wzi�z/��5�8�;��$�� $����@��O���ǳr��Wo�+Blxa������v���f3L�tb��Ͷ��$�����E���4	C�(���]����u�V��eP@�,P�c���&Q'76zMXgd��k]�S��@�>�U*��ܾ�G?�U1�:o5]~3=4h{�}�k�R=�2N�\>s�WC|��m}�
��
� �=��l��#��f2��q��fYp�J�H�l�a(�r;�&/(�G�5#���x+�06m�:!�05�s�88����N�(�:��p���:��� a�$�L##^��F4D��>�њĠ�MV�/�^G+*%�)�4C�o���Y}���<�F?�U�K�6�Xse ����ڜ����TNYf+Ȓ���l��[n�,(�F�&^�l�� �Y[�J����6w��?�(wR��jt���o�q(#`����|��?9��� o���7?�]\�d�r����<�_�6�S/���>B16=�Qߝo�^�Ŷ��h�9�(!����9�Q#T�5$�"�U�,���˜���#k��M�o�^�N�FzT�bm I���Փ�n��p���Cm�f���G1XC5H�r��y�-R��Ȅj�A�P�8|*��랖�P�Yrv��ƞ�v�,��tɆ̈́�@�n{��V�G�rd�����Y������Z��m�����"��:�Z�15*K'(Э�҉�|������г�Q�sQ�n] ~����X��V<uč�%�D�q83rH��2��APb��ƌbn|�k.-@���rR�r�Lž[�?�m�K�8@��x�V}��F��Ge'������Rb=[�Y��jb�DG����)�AG�5P"x�~o_�e��R��N5x��k\���S �[!o(���D�H�yV�w~�#O��邆��cp�GhV<��w�J��c��ʝNq�(W~�)��<�~��v��x萁�\�Ln��m�9����vG$E��
�`!���Z�����'{���$SU�������X��������� "�n*C{	#�كFI�O���<w����vZ��߹����+h��gGnL���{R���<&G=N�<sa�0�ƣLy
���Ӳ)n�.�)�R�!9�r�5^v��^XV!��1_�$�՚?��4�
������)��=D˃	ʾ�-?C�iq@/�F:����4�pj_G�'�c���ɡ��BIJ,�1�b���[/(���	_c.qK�)����X;��K�� ����,F�+�{�[t�ڪ*�̶�<Kǒ��I.jlq)fU����ϟX�\G�y����5�4��d�%*y�i���zel N�Ƃ�p�)纱V�:��xN���@62qU���+���C��n�5�UX��۾��,x|l�&R�-���4�Np� �x�&�����z'�S;0g�P[궁R���(I����;7 ]�a?�%�1�$�8� >C���T�6.D�v<��U`Hr�?��z�>�(���6`v?w��>�Z��(���pu
T�R���W0�$��h�&@�os�	Z�&��@ͺ��i[� ��<n	�v��B̤��z�M�����, �4U�5|ڂ�v�C��p{X��/r�^��ϰ����풙�z����XI�DV���sk�_����a�{9���9�ǅ<����f��?���.
<��:�ld��1�v�W��q�2���a$u��Ӂy�(X@F��uq}���cd���,�D��K���Q���A��.म��
-@� ���}_��%X�I�L�.� �ǆ~R��Ꮕ�"آF��0�w�Xw5M8��j�"�m0Q�Ό��ws�dG�$$�:����ʏAu�	������r�L��%8�b�ͫ��#$hҴR��MþѸ¿�P�F�sEewñ�*}:?��+��D�ߒD'�q��eٟ������l�7k��;��c��a37�҉�*�2J��>��$[��hC㷞���@)/�7�`A)��P������4�:(�"
�J�\[ &�x)b]���x�7
7���Hn��}�<B2�B��2n��E��<ɐ�
w����=����	v�H˽$'�))�WYՂ
9a&�IR�"CD5�I����H��҃_�H%��e�7G�� �ө�5�sd��O�O7�AH,�s����Q����^���(�oG���b�����$	˺A:0��� SO�N��"���㔲����Z��
{�0�m�0���@ZaO��0r?�Ơ�����v�%X�@3�8LCT���+��� ur�!t���\&��{F����Ht.1�5*��d�l`eΑ�F��G~e�ũb�W�zw��&��B��o�Q,$�
�x#��,Kִ��d8V[KЗ������?�YkKwHF�g:´xv�9B����I��*��6��YG���c���ȵ��r�"h�G�CC�CbhR����?h���R�q3�<���+N�u��t Ry�+=1���7�B@A"�w���Z�|���IeL�x�����>CS<'O���a;��bY1�����"�
�E��6x���?������낼
VX��s>��w -Q̰Z,ѧQ�A��Z�����	!��oh�:ğ�7�a��۟�J<n9����:7R:��Y��HFK�O�I�	���$k���Q�Vgq����ɯ�,�p;�R�c��B�����B��:�!�u��՟�nv��t����ȄݡN��:W+'��y.�X��ɊD��=F���ߦ���Vk���x��#"����3k�T�f?�V��xj���#��:WB���P�)�7ψN
a(�|��(�@��s��sR����"��^{�`{ׄ=L@�'�H�N�*]��֌UB�uBjIК@��M|'�W]�E��=�3F�+�X�!@�A�@�d��R�j[^��n��kfV �$Q^G�����`��ǫ�$8Z�	������XI�G�i�U��>_�d����r�}1�5��`��m"(�乨_1��)9V�K0)JSs@���*�)�1�]G낉���s�M�:��f��n�_H/=�Pa�Wǜj�4��'ǵED�(��n}�=��C~�� Vz���'�GQ����[�J*���>Cm���Pʦ`�gj��D.�_�:��*iU��P��U+��Y@bMd�}��O&�h�w����#7\����(����nq0b��I��UK�<A4� ���<۳=R��տ�
�*��ZP��Gp��%@�I	��]�E�v����m9���T񢸁�p>�F<�
�.k��P�E����t��Q��hP�k��d�^31���Ġ�?�G����4 �@	��c�xs��|�x����lJoț�f��) 6-&�;:��0�3�$���r�Z8u�k��T���8,�BA�R�:m��.^g�U��6�P�3���]���ǐ|M�g�چ�fj�[�Gh22�
,dU�iz��t'4Dupk/)�j�o�;�*B��O����#���Y� �*�]�C~M�r�x��:��r�;���im�y�5����a70JY�b��p����c;?6��l�F_է��l7	�k�'Lx����ď�TM�3��N����u��F�� o�-�	�s�������4�Nu5=�Sn�t���!��\nt���?�/�W�5��X�g�R-�q�Gj��4}�� S��6�mp���ȝ[B]⏻�-��p6�����S�5)xVQ�� ������}�����}�]tc����K�V�OaZ���3�z$nG��č�h}(w�.�0�
��~	����D(�ā��U���7�&�N�p[1��P��	-
[oOl��L�?���.��"*��ˋ�C~%����B�UN]�eפ���x�L���x3�6`I�^��q�,'�;Ji�BDJ�����Jt��NK	�����`�[5i!~:l��;�d�Ek�����T��WcR�7h�,?�����pA-WO#:��Z���K=��`��x
��RO�W�w\aB�\����7�I��wE~v�0�J`l�ר>U���G�9�<���o.�����V"P����47��*��`��M�c�^�5%���ό����I�t�	ȯ���k|�RH��L\3��pkC*�
��>��;�$���o�8?*��	�6���l[���	�=לQC
b��Q�� ,y�C�1=��J)I�a�&]���x�s�)��M�`?$��AOs~���53p�,`� ��Yf���^�wY㯾*1����#H78;Е�8���>��R�C/?3��H��pp����	4[e�R��TJ�qMd"��a,Nι��*jhz>����&^>��Y����VR" au��5��:� �}��x�����z��/*T��D�bo�5[#ҍ�� ����[��6Nk֡&FK'�Q!�jද��Hs�
/R��[%��o,5��e�癜�'2Ժd�W0߸�gj�s��,���f9�����\n��2y+ ��-���S�v�]x⛽�ƿ,�U�?�����C@�U~�3pM���3�I%��gK�D�e�\��%�ւz�/��ksvD��,U�+l?�1]6�)HP�P�����.ͭ�6J�1���7@�2s���t�u��F2��O�](�x�.%W$T5�i°�k��V{CdUc�Tt�(˳)�8N\�@9�2�H�a�G��&.E�A�y�)\)%c�hLX ��|vS
��F1G֩���t����B�#�G�;
��J>L�7�\p�ĝ�J4-�RPoa���ne{� ��'�O^ES<3�?qi�O��z LzCr��-{ы�/��),�B)�F��q�������s�Q������h�wHa����c��@��=+Y��خ"F31�ˊ��3xk�h�o�!:�W����~�y�p�^��J��Ңk�)ށhuc�՗ȳS��� �zT���)��o��`qx�����bR鱤�V����j
8V$1>=��Qx����N�7��G�=��ץ����I������CY���ˤ�c��Xgv���~��M�ݡn0�=N��P��G�ڻu.ȇ�R�-�i��m�nfu�K��¥!a4��s��Oz���$ ��?ߘNdۭh�fTɹ��9�]��0�\s.����E�P������	�$d�"�V��EK �n�.�g�t���C�ȥϤ���O�Y(�;�5.x�|y��x�B��_�r�����6?�`�R㼧 l�m��Ǜc��vQ���n���>�/4�o_~J0 ��
��[�.C8�cw
�0Zѝ1��r
E	�:#���AҜ��j l76����/��+�/�3�hօu ����	nu�x��T*��MN�>	/��>�G��$��)<�#�Hj��>��T7L�z��l6>Z�5�����2��i�uϳF�� ������QY{_�����Q���j6ߩ���٠	�d�9�6�G(���^��6gd������y�2��-��Mp.2�����,��w�-���ҍ�E��s�	�6���ގ��#)�W�I�E>��1��Q�C(`l-������y�ףr�c<jku��?�ݍ={6���W�/Bd6�P�7�,��H�6!����O�V�p�6����r=�&
��}WFCQf�]�$'��-qNSu��N$���E�"h�G](k�+/����dj�3u�c��m�*/WF�@��h���5�C���4�.-���>^Kr�́�H�Ո��ɷ�ш�$8�lL|֙���a����y{~e;'��>�t}�I�U�:��/����bD��ĺ�V�]C��/�NЫ|�&���(����\F�ZBi�K�}M��Q/�R��IKsM!' ;��h��V�ז�	��Q1@��c"0���֭J�#-��$?��#�� "K/�O�"9[?W������Ui��4���(����������^���/o���@��d�0-{���O�wF���%�}�H�N#W)����\H�5�m�Hc18��=�)�����G8��5 ���!�$�c��P�~��ɸ���=��1�U�=��N���4����
�{}p�jq�y��8�1^�j3<1[�����X���N���xl�K�rP����
ǯ��g��%��	h0'���o7\X��bN��f���˰�:9�]�����Oʏ�kF��|#R�+�V���������έeF��(YU��g����UE�� e�3������&&� ���%���eo����P�w�P�zpM�b ����4�MS���-U4�@��/��.R�D+��4X
}`���)IAL����,Ys����%��eܦ��F��y�qIR��t&��HeI�5��2������68���ʧ��J���oA�[i�h���KF���R2�͘*ԥ�;�0�<����)�S!7�܎�T�ˠ�P�4�������d�=o/~ �܄�@J<{��J�P�v��`]�z�Ѿn�|\�2�U���s�w�Q��ߐ�F��w�A��s�T�w�<�	�J1�l�ą����"?��d+�F>��/P�хx�\��@�0-����[G0�˯�ё4�6�b�����h\,���LB&i�y$k�,v���ŐGrk/�k�Z�{�y�N[Q?�vpv�����$\S�Ip�B0Қ�gތ�/Z�v;Ӗ����$Ʊ��5�Yu�D���H�j�L�'�	E�5�������	"�)���Pp�x���^�lW4�Vr˳eS�d��ny���#���W	9��k1�õ�j
^������k���C�_I��g��<�����	���� Ԁ{�����bIo�'����dn�o���9�t��2��+�!q��-נ�����ғd&�G��J~ϛƸy�r��?+�z%e�,#����C��.�J�cv-Mِ�7���IAE�d(R8W1Vd!�e�������Bhl�����;D������_��g�	����!��������b�ђ�4@�e���Z.GP�)A]_��#4����z�6�:cN1nMy� ��{F����E�b#r�����5�{�B�w�:�1�/�n��mG��'h)�v0A���;I�[�6^�04;x<e�k����R��za�c{�;�"�:"g��e׆X�^H�Ul�Y���L]|xѠn��>~	o|�f����ӿ�lؒᴧ�K��5�E�n�߰:#bڣ��H�7�>.0Q��ƅ�
��XՏ9��f+���\Q�nrQv�m�b������{K�sk�~AH@������Pt`�n�-p���]�p9)�ۏli�t!�K�A��G��1�i�Jp�h����*=���y_�!)ߙ>�`�^)�F��r��KH®S\������P��`_f��)ZW�@�#Ⱥњ��r�e��i���,HT��j���IM��狼hXX��x��wSx�-�&��Rj�~�@�l�6��0*��؊z~�Fy�ĥ���)�-����p��pGo�p$_��@��,O���8^�[�4��G}���a�c�5�
�r喞|��i;=�eհԞ1e��Y�(i�jt-�s�h}�|�43�Jc/���n
�j��g�ӄY�w��B�'%z�^�#�`����$�R�ͭ�"�
M.��/c�F`8��c{�>�?�����Io�����,�gF�Z���/e�=Is=i��MzC۞=����¶O��j�sϣ���߅��Z!ߗH�"�̽g���h���f+��J�.�=��O;Ă(f]��Ts�'%&�F��ĿM��6��)]X�r����pOAa�z~i���GDw��wj1�m����ԑ�w�J��F�5l~C��S����A�WLp�x2���C�'Et�*��W�t6�,FR	��/���_���yH�c745?cSM�t�o�{��]�QGD�~��)L�
�� �fF�VE�pr���v�_���B�$��P��ڶs�����0-s���Y�q�;�K�)���ZHNX��5�S���sm���΋{��G�v�C�2����)R|�7���nD���@Z��jՐ������gZ����M�&���}wQ�L�W�c�F�Y~ޞQ���5� lC1����?0Q>i9w�bl�a���[,��<�!���ɼ_��so����t@?V�²70n_�7���J���])���Ȼ��* _)K�cDes|.|��rʴ\�.gu,�{��5Z�w�2��W1�^[Γk��5v�����(���	m?�
O|�dƱ3����L)�b�@�m�,9^X+:;��gO��ӿ�u�u~z]��ޯ�G�a���ȗ��nw�V�]��ZnA�-n����BB~5�����=��Q�������_�`�"	�"����,�톶��x}U�����o}�D�%v\�M%ty��B`H��|���$���_r�Y9ɻ�3����՘Xc舘a��/����oU�ڪ�;?��mp�dPJ-ؠ���V����{l���\�-�Rc\���;Iu3�����@��6Y�hL�u8X}��rL�<љ���g���^c�������=�niiem��W�2�Mi�	]W.�ts��W�&�GvD{l���>�+1��.�)�M���K�k���]ܐ�!�\�j�|�V�_<a��IP�ԈY,�����XQ����`�kR=�	�`C��xD�/=�I7�nz:�����@�>ۻ��=u��y�w���
��*sT���UL$W��H��W�R��
��I�(�):���O=�mC2|xf��5�x�D t$�3��:�/�O�	�4,�Qh&? P\���1!g��yn��hf���kue�J�S���8_�|�ͣ=��cb�N>	��S4V����{p�p�PN����tX���כ�rd���|��I�"t�7�M�J��5�9y�p�+��6�z���t���v�#4��[]3���qs���k�t�=�4n����%r�D|��fV������Z`ŋ����}5'��bЬ�\+�s`��"��[�h�� � �2l y���8�@��L̽��i�����̿��x,�PЫ�?b3L^�%Ļ s�;Ш�V%��]�^��&��OY�hi��h�,�hmc�1ú8<��pYO�*�P�[�y*���U4ώ�}����t�ߘA���[��������!םƩ���e���S�D��F���V����
��F�K�lu�q7��2��+��"z����9T���<I�=.*S� �9��h��i��Go:�t ����8�E����~�v9���a铐����~�]�B(�40A[r��#����Ux��[����v�z��Jב�`�ee���:B"ԃ
���_D�ה
?�c|��^V��Vr���=L���RP�T������f_Eyx��¡i ��~r��-�;g�0g�5�Q��1����(ܓM���ԓ"��R13������Gt!�jS�������-%Q����Zک�]�G�Z)����?D���Hm���-wm1;��q�L�����Y��6/�eܾ��t4���j-(<V��Gr� 3��e@����X-O4b���	�BL�B�_��қ��	]���~Jt�:����KC�z�ꏛ���>���dy��>�;�6���[ҡ].&��9�9�[P�4r��f9�z���*h�a?�1$
���0�T_�	&����=��ߌ����u^� �N(�+@���h�-V�d1/B���(F��Q���[��f�gt�Ӗ<�dQbg�w��|9aD����[�6_���;Gz
d���A���.��x�g��5�
�m��l91gb��]�E)�n���(����n8d�fĄLv]*�_�E�$eݣw�پ�o��3��Zz#����j��b����~C��}'�,N��_��5�J�kR�_��N-��Q� �Ih�� ����s����g��o��rtR�8�]=��`�55�U���d��0�_W��i��/�:Z�9^�^�`.P*tx)�.�����o�E�=��WYn��I�w���8�P��$��/����M��9
�K/�V�'��0ͦg:��Q���4:Z��.9e_6æ��[s�����e��A�*lG�g��~Z� �瀣�'y����e���X�������KQ�Rߨ˖�V���'[v�PV&�@+���sr�$�+�X���8�x� n6�'+�[�.������t������5^��6J�b|�#(�	��WX��_�>��*|D��S���~>x��v⹜�I�eIFGRQ��+|�9�h�}o��HZjtFHG��(is�ܷ�c30o��G�]�s��"y�'�%��S�Y2��1��/ �1��)�E�i�?Zp��|�ÕCr�Y�Z��)�ω��gW��lf���@�<ce!��ѧ͊�yO
����m��f�#x�Dx#�ttD�4b�u�v4�����%��A�rz�Z�3\&<	���2��*":_/[�$)j�N�yP}k�����T��l
����<�
�%P"z�W�.�a=kQ��,���FB)M���̆����vv!a�Uάq����UO#,���i(v�z_�F��]Qj��PSd?���KՐ'	� fc_�I|)D(j[C~���� #��v���bJ<�[�dO���'D�i�Fp$�0�5�ϻv��0��Ҽ\��QX>�/䑘Ŏ�i�}��P�8�0A��\�����4d-�I|:�l����T^����<�3�?/��Y�S-3ȴ���0�]Ü��_�,d�U�6x)y0�㛈��!\v���c׭��ƆhqP����L��Z�ѷ��>�<PR^ZΝm˷��������Zq���r,_o9�b����[}�w�}�Y���P�\R{�L�%{�y�#�1��dk��W�;U8�f��/�C<o����*��J�;�b��o!eጮn`��י�ԋI����]���T%����N.��k�Fk��:���Y)a����86S�{ʸ�9����G������i�bc�'�z�����n���b�l���4eMM�I𘀄3�����͎�h�Wʠüϔ���G�w��G�}4�T�{��u H��ط������;ܵ�OY�zo�aɂ9��a���=ho��&�A��k�|�x��-|�oy�H(b���:������zo؜Bc�!�I�c��MZ�\ۿ�\:q2�*=ԁ6�w��t9���k�د%^��Pۤ'g�r�Ŵ@��Y��Zb<GÈ���+^q�T�ɗ��7����
�w�~�P��LҰoc�J�~��m�*<cER��6��ϙݞ1�[��D0=���ʓ�r��Ǘ���`��=Lӥ��yO��̰	X�-��~A��4�-��7n�4t?�c�χ>�&Y��[�[p7�3:0�ߓ|�IWM2V���������Q஻�1�2-zlG>���a�"k�y'3��:ٞ�E���?>�3ryA΂���
�H���v���[kl`\o��2�2V~��h4w��F¹I�bO��L`9�rhI�ių*\Q-,�� �
V��[�������<�m}�ig�PN�cܧ��b\XO����o�j\��w`�
�WIm=�R*k^D�/7����T�W���A9/�����}+s ܙF�n�۩�'��2�:s��kԪ��]��Ӷ?JC��q�4��&��M�Ri��]cW�U�H�n����X?���Ο�:\h��*SB�H�ܜ��0BZ<߯��#����3���49"�;#�q���1\$S�I�a�E��eC�������h8�j�]�؏�&�%��
�S�gȞ���>q�n=ѽ8w��M��h��kR�o�ZWPi�t�K��Pp�� ,�Ώ��	��@`��-$���5Cn-�et�nl��8�>�S��������)��	��̸d?+߻[���j˛udgX;�/��?�VH�K�k��\��6� ��mv�V�C��.ȵ��C{������o��m?���7t
"�&����|�C�V����.����^���*#��O1��$C�2���y��p�M&8�_;�P�n�����<�t$�h���{��xtW�P����f~�ܬ~b� y:\1�[��7w):�n��ɖY��㎸ B6��Ԭ��{�Σ���+<���b��ϔ��'X����EH��t�@N5���`�{3�
�L/��?.��$�J��ؼ��5���A|��0*��@���-� !��6��XD�̡»��D�����@�$���̀0���Zy
8�3)���+��.Ꮅ�>��$��$����O&uE�\� Lz���R��o���6{K-Ny���9��t�|a;��N��i�ho�9�f��5�凶c�!�:��0�v@�׆���@\� �M��Y8cO�~��/q�#k�z5��X�G���e���UO,�B�2I>o���6d�4�k�Usۙ��&�}J���ޜ&lXi�'#9+�}��`!��S(�:pTF�x���헇޾,�=f��ky�h�����@����q>�Q�L��`3U1FM@s��nx�F��L%g�m�:����9�J�{]W�&Bw���+�g�#���b[�������Q�����9r���S�?�9�U,w�,V����t�AE80`�`��/!3�q�F�/��)
�̓
�RתSf�,ܗ#�+G�R�FG����@Q���N7�
b�x_���>-����ទb<�'Ϡ�;n쇦�E w#���ہ<�f�5����َ�P'���g ǃ����]��ңρ�q{�Wыb��_�L s�Z��sT���&�z׬��S�== H�џ�'q����m{�g�)�]�{k�e�M5��33��\����c�j�Բ���f�$����Y&�$�uRL�R��$��tZpD-o�y�� �k�Z���Ԏ?z�>H��T�b��Eד�"!��%���ѐOp@b��]!��T+a�?X�㜠&k��9|�.�s�l͘5f�7�(�ƳJ������ɻ�XkV��o+E,T�¤��pY��#�؊��1K�[őm3BɈ�;��Y_�w��{�N���M5[��W&0�I�3�F�]!�X̬�Ǎ��P~:�)� *_�	4�.��X����ꮶ�vFb SQ��>�[���l��U)cz�^$�.��+Vl�����V[�B#r��0��Ÿ�ޑ����4�I҅����q�0Hlƭ�B�0A�M��D�4��չ��@E�J���u`[�U�Z��/[�׈�����I�f���xȠi���G`���Hf�!#���<y�K�lyh�r�-�f<���^eDkٯ���dwu#���(S<���� ZFjJ}�a�ڐ�Y���A0����:�^�
hYt��)��a���vR�n��*o\�w���dC�y�+Ҙt[Ps�OȜ��X���!�r1f���j��P,|����e&��UP.ڴ8�#?A���'�݉�.x;��G>�����!a�HRP�����8;�&Q�%i�We:�;1���u��8D��l�y9�����ɼ��YH��zH��c�{��;+���s�Z5��|��2�t��Ru(�؍���̃�N�r �H��@/��d��e���k����,�+����ëz��v�u���2���U�\;�s/�̽~�oT�zr�e�[����n���R°���*��)o�Zt~���2=>�8
'n�:I�n�q�!~�T���8Rn�m��#�\ˤv�)z4�]��bv�s�Y?�v��Ȏ�t$���"�gC�E2o���@�Qf-i��{ڑ4�_uw�4�������F�p�*��.��3$�+�\�_�z��������s҄i���������d��-��|���} ����
�J�-��X:`��a]�5.�q#v'T�c���r��lhq���)��(|���P���j]ɀ�N��o��mgxKWQ���G�d·l*�����S�z�TDŽ�x���Wyf��*��)C�DOPr�.��\WTh��?׻������/H��7����MR7?z�3�u�Z��ѻ��k�s T_��)�.
X]��Cq/��9��<೩����o���
�%s���K®�.s-ţխ	�Yi-�1<T�
m�Y"9g#C��#�6Z� �󶽴a�Ɯm�$����{�r���U5�G�
��b��<�}4�>v���"!7��;�jh�W�ѵ8Y�/Z�5NW����I����b=���+�Q�d���E�"�, �c���I���)��]��3Eg��8g���֕���X�i���~��zQ�z�N���=j��*��^���V�<�Ej}�;|sJ ��~��J��Řn<����}��_=��f
&`'J�l��0���-��tۋ��~d�?F��i�#�\~8���ed#c.�tT�>��r<�ca��O�Xw�)vB�S�j)��l>^�ڵ�أ,�(b��������O�0��=�����#�|���,�������4M�qr�������u��a�=T��L��^|��	���fvm��]7z0%a���c]�2� :��M(��b�6�6%��\?G�M�vv�P���R���(&^W���>�Af�N���fc�
1��@���K�/���{L@ �����}�j��|��@_P\��k�hʳd��\��ݢ<%W���o-�Cm���	�R��#��+��XȄ^*�<�S�I#Y(�����3�o�ޣ��pE��r=
�����`g'��*�/��VE�/D��!��#��5Yp^�F1�P����T����I���߹�&@���E�<�)k!<KH����z������	n����G͑c�:�a
Fu���3�e���\zu�Ѧ`��Z������?n���x�����.\��LF�|��N�H�Q!*�*%�}����B�Ң��;Hw@Nݺ�������G�q ��oBb3�>W�Hv���14k�hG���7H���	y�`�Tŷ��J���9��\�z�:���Z�4.[i������ݸ�ڷq�+^�=`V|{M��S�(-ݖ�3����%�z:�9.<�VV��/��%���7�5JI(¯ۚG���c��8��g�<��}|�L���mɍ�+°�#{�/MtI�4�����U��ޛԲ`���c�b�$+����=�������h�b��X=���\�ނ���z�8��[��X����G�/�D�n�S�����>�G��P����vr�d'/���a��a� ����DYF�Mp��o!���6-�
��`�6D7�/Ꮸ��_��F�݋��e4S�fK�]"�R
`�p*���jphW�`�6�q���|� ���9��T�i?a/:�)EGz�R���$~z��!(pW{
j�05
m��I��7�/�TXHX��Gb}�j2za����ױ�G�ؾI�-�����57h���٘�o�t%%��N�	
`5OF?؃�/�VP\T�7����Gk���Rz6�g�o�l��g�����ѡv(j_�˧��nP7�(AO��f� M��p7ׅf��
h�!�b�����ў�1��b29��ł[tb!"����j,���Ec!����)}i��r���Ⴑ�e.	�a���{�钢��*{tS���?Ppf��md�c��u��~����X. F�S/K�3I����
8A���Tև�5��~Q��_g�v�}l���F�Xs���
�����@�� 9�?�PQM���3��
�S�,' �y썌����.0��#
���~!0@�<�D:�g�u<������e5!�ƎR�Oq��7�v�o�.���T�!m���H,/�&�C��ͿM'�#��HeP^Dc����H�n����?� 9GK*y�q���6BQZ��/���w p�z���1�~���#��� �����Tv�*��o���S����X��Uv���Pl ���:�&'�+�l��1��}�b��u�EG�GHg��x��@mhD�Xk�Zd���Ҭ31s,='�G�_$�a���d}�o�H�(���c~%���2�h�����Gs֘݉>���V���x<�����e��!���j���ȓ��^���$���$����
=~���n�澆x�	B�(Dձ����6�؝*�̿:K�J�:�i�,H�)�XBO $��a�i���]"��^��������-\��Q��I�.�A)Ă�.\F���"�ߦ�3f��X�J�*h�O�Ld��]N�p�¶�k?�@��>U��9�YY���o6MYqc||!#��"�T�8��QxT�E�.�FH\FWQr^[A	2\u����o����Y�L�����)���e��F�q�[���� l�\�>-Rp2�^|Xl��K� �l���'�I.A,����=;�G�)�,ʏA:h]�,q��Q[v?Scrs+b���w�� @j���l���j.��>��[O� �
�]�8*bU���*��u�0�e���ާ��c���w�F��<#6�;C6!�F�ŉ�J(�I��;j�9K���aβ �t�7bl\�Ֆ���\�X�94X*��I���|�e0�W|w�\�ʎ�OS�Y��jZ��H]�G�`�jW�V�;�s��GR���giT�9i��X|��<����C�6����i�q�bx��3���E��u�z¬��3��Z�ȗ�4�(��H�݀��\�����qy��6	b�� v *_k��V��f[E1P���1u/2b�,��y��'|�a ��c#كӽ��u'�E���ʀ!O�P$  o�)qe�;9v�Y��ƒuJ�"��=�k~���ӐEA
:�v ���M7'=�t��;^
��h*S4gsKۼ��H~�v�D�Ѿ���[�3bv�l����*e�^B��ˑd�\�����Dk�l�V�XB����w�}�*��M{�z1-$C[FEtq�OB����d8
Ș	"�}��ve;w��sG��]Vx謂���<ğT����P~�R����p���H�i���J�l�T<�Y+75F�K��m��-����[%a�բ�'�4��bj\K#O]ى�xN#���ڪ����#ٞ=�4fD�ů$Rlq�4pvh�jv�ZJ"qS��� ���3����n�B�֘;jvz_��.y-�}��
�N�x�J��?[�ڶ'�6�_��9Ӊ�/>a�9���
�݊_��9������a�hݨ�\8�+��|���U!{��t��D�k_��ʎ��}��B����v�yA��l��Qv�2(�/G�`��浔.�6���[��_R�a}լ>#N��ѽ�$x�b����y�f�
@�%à�EĊ�;�x;�
4������j�y�{b6����*0 ����[dB�����{�a��T�ڳ@J5k��z���m�x��px+���ڜ���5��4S��*���KP��)�h~��H��[a㩡�jY�i�l��n�-{�<�<q��U�g��' !��ʠ�L��c��V�����T��d��#���H�d��=5���/�%�3fF�6LZ��2�G8R�$����V����:��U����&_�����8�c��᭜����w&?�%J���&!fҷ���=���r�]�ҟ��M�H����d������f�&���A����~~=j}��W����$0�j�~�E����^W�mw`�O&�ey��|h�qQaB�7|V��mj�)�.�F�	˙���g�N�\�.����^[�"�)�sH�"����ˏ=��t�#RVSz�$���wγ4[�m︿������YUL�i���'� ={	�R��~ɠZ�eb��ɣD�c�0&r����֎d�����]	���R����ܢ�Q�\�d�i#MX$8��4;h)���pISS[N^H�j���sVo��Ix����Y�k4�Z��Th?z�p��B��ʲ?���+]q��/`kb�ѭ��4ڭ����$�)+��۪5��12.�BS�����L��4<�U�߂�9I��g-㷦�̋��F S�����O��/3K�d\7��Yp�A�����L־��<��� U[�(�T<|��m"e5`շ������:aEy������Q��BA+���#����}m�Ӆ��bݦ�4 M�9���P�&A��T\�X�b�i�Z�?����J���@AC�D:<�Ԗ��U��.Xm��p"�"~dH[���B�����9Zl��A�y>��b��o �L�$aԡvc,��tɴ+2e�rHV�5&�	��O+0��%��`WSb).��:�<�j��QǰdnЄ���[fv�a��L ���>���Qq�Ob�3��(��ьb�%+�n{
�BÉV<�@��" M����nԐ�ށ�΂�(���e�X6�N���hBv%�%�Ǻ�A3�D�8	��١U�ۮ��N �i~��O>N��];�qkh����eXӧYz����ز���.ܐ�q���"�ک�����0��P��s"k<��an� ���;0����1
k=�yJ�6u��/c��Z�@�
���(��n���4
�C+2���N�O��X�E�(�p�;���"�/_���?���`h�l�-�J��|��-�kP��b�3��'�׶P��}N������b7O��2'g(��6zs*��ˆ�1/SFA�d�K�HN234 ��dp\�����-6�T~3�������ׄX:��!K�TW��}8�N|��Ɲ��r���6�Da�RU�ig7���-�7q��w�f�U��Q�>�)���;�{lHA�Z�OT����a@�~Z�woFݽ�v->�N��[qS	���	�<c�� �f<F �k�\�'�*�г��$���$�<����1E"��~)"l��iϋ�Z*�ǜ�'0 K���Z�X��μ�Ly��W^�[&��"�@O����م����������`�88���tf�$��Y��*��æ�ߩbmX�0�T&���Ól���>����*0"\y�9GE9h�<�-f��N���\CA���"�g�����qӚ߼c���+�B��-���;[=�e$c T3�-"�->�ܐ6T�Q�;e�"�Vb����*z��4_
ϵ� X;��\67����t�~�4=FY��Sh�������xf����a�ne@T�E'��u�Kg�}Q��>�=�8׭qS��8�n9}���i��ԭ���N��%�B��]{j�FKmϓo��"�8a�$�^]]p-Ä+�����qŢD[?��wK�F�b��~��(I�"�yF�r6:S&�>#
JiY۰������R�%�h��i��k�X�|�:D�P]�O�^�S[r�pF\�4�"�P@zЋi�����.���x+�p�EJe!��p�&Pգ�Uܨ�%��A���� l�*j 6�jJ?cRw ��bnUuȪOwXإ}�%��j)���t(DT�tH����7�hx2����������C=�Ƴ�C�7�~ݖ����\�3ڑ6T��+z�����I���+g����8W���L�ئ�����`s�W`�T��lSLܵyҥ���(�V�����N��4�CFjوNw��ޯp��2��E�o���ꓬ[��Ru���� 4[!���չ�o��&�s>KW7���\E�3�i����K�^�Z	��`���1a牣h<,ʊ��C�,�JH��'XigxJ�w)���v���w�N]+/��ikfU��&У:����i`���n��+L_���>�e���j������u��~^I�:=�Tk�(���{�?~�wc�����J�%�ˀ�����Y��Q����v1�BI�{����<e��b
�x���'���c��9+E߯�f!Ӯ�k���bG*\����6�z0��xȤ��Z�0���&�U�g�٠<�b3� ��rh�K��GGu���.���И��y�yNu���|�af����8��S���A��u45��OS+K�U�I�k;�%��x��Hۛ|�@��y�e����Ak���(��oY(gzia;�]�[c����������=�@ ���[�u�碎��^��k���	_I_�uj���:�i�_����X��J:�=�e=�ZW.�{�K5d����JKX>�R>C� �bo_��'=�T��)=�͒���h����ͫ�m m�>�и�]$���{�Ғ��Nri=k����aɮ�5aS��$<�����."Iϧ���Jz*���pn�}�QIٟ�~�϶N�ܧ!���l�tC���� ����@�U3a�>��A�8��fO���4��q,���}�8���>�+u/'���%����2����ݱI���|w�HP��ٸ���`<�x�o=��R��Y���
��y�][��򊃧�]��?���Eզ�&�(�T��x5�^7�6�d�D��}��kڽ��o�&_H�@ b��2D=�B]Ź8/�h&�l�N\�����g�}�.�7���v�m卭ג������aT��Y�DF�1�����=9��]�ÜL����E�F��4H?������H0�m%(�V�wxIK'ؗcF����s�_^�?����}z!x��Ip��B���*@m�z�2!����#�_���B����]ˣRğ��}�ۊ��mfl��{;���U��X�j��Wl/ >'^���A�8�s��I��yv�ܓ��\O���:۰v\�s;���=�K%2{�c���7NT��zB�_m�����j'�3o�vMLf�~�L�h+�T4�MSc��$3Ҹ~�Kl���ƧT�x�C/�q��`ߣ�X�Bl:y�I�	��$�f����K�`�i%1.D,��Yn{��̑�gU\6�|���8����kE�JM�A���=Ǧh����2��ó{�f��2>��
��>�a���k8�Mם�yL26�_�LΘNr��gQ���d�_��	J�).�j+�a��}�Ӛ ��eͣ�TُZ=r�"�(��,>������)���\�1�T��K8�h�����\���a#��IU2G/�@c���7lJ�=>ځ�!|L71�C���6�AA:	�<o�U��I�j}�8����X1��ά�Vz����L��m��\������N&`�ؑ�Q�~��X��a���K����4I��:K���B�̘�~}ѢL�� O(_l�`�tse�K���o2:yFN|2�
>������t�B6�����P$(w�L��Q�h��ݐ�b��@�����ȱQ�y�J�R�4˒�J�|C���O��j ;#-��u�ǈ�,,���P6�[y,��b�,E���dQ�ȑ�"}��q�ւ����q��OF�/�Z�5'b�]���q$e+MFJ�ӳ+y����9��l����D
�o+oj8�9z^��$9X��By!)�ݖ|�j�H�Z��A�PTNoU4��*0��/�&��ڟ]�Ms8�Q��+��5a�T���� ��]��>�B3=3�P�\H�]��o��q������x� +�#���g��"���/�R�/�J��]z#&�O|�4�i�Nk��!	(6Y��>�ח�=��9X��zͷ�{�;�ŋ7po�l|Aa�ɉ��#k�ſ�c9RS�K�F�b����@m�7x�sh�ȥ�B'oWC؃T�Bes��ob�ip�*�+-"z�?�(:�L�Qm[��Y�Ud�/�m�ŭ�=+�O�Cx~`Rsb�����'�)��$\\k�͘�����H,�-�7pJ~	����GPJ���;w�p�ݏ� ��åHt�;�]-׉E�طz$��
"A�ю3^���=�a�k�r{U���!Fj1�����C�i)T|H�WT�SS��wPf�lH��= �0<~gJ�h��$d�u�E����.�	"'�JF��,���<�cJ9L��A�2��vD�Ƽ�W!���
L�������k�Я2�x��\�C�W�u�e���続�.�O);F��r��0�$15g�,�Ӭ3��f�I��ə ���xbNP��ْQY򅔊�D�� ��5���*7rU0�"7�Yϋ���8�v�'��ngg�bG�O��S��Z�����h7�O@�)�W5`��̤��B��l���D���Q'@ �0�t�=v�Z�/�T5k��s.��sHT(����~�Z���I�f���9���|������a����*��oU��A-���m��yj��Q�?=W�my��GK5�#�O
�|��y4�/W��Xҙ�@ZY�xJhq&2s˦��w�腀gl�y�Q�8�f�,����ע8�^}�5*�m�8p�uI�(&�#�-���>Rk"	 �
)������e��+I�C�r���
��Z���A�^�\T1�
�M��fc�&*�Ց�T�Q�:�����p Q��lE��p���6ƪ36��y �ѯ�7�[jf_�ɚPp&�»V'��en]�d��3�����Z�E\���Ke�
Th��\H��z�#"�J`r��$<:�㹽s��+�o�:��y�� �e��2�L)DA�C��ġZ�" Y<�;�C!�
�6҂(b�A<�*��_ㅆ���ڻ u?x�ܤ2�, ���P��w ��B��4�0�j�����6�
VO��8h�ʦJ���^�J)�d���IU��w��0R���x	��e2�:	K�;,��97vZ�(���9d�$�ǤVXW��T�I��E��ÕF!8�E��P���l{LH<:��(��C�����,�I�
������_�R[!θ��5�GkS�Fa�'��\�\|Ԅ��B������7�����ɽ� ��,s�IY���w,C�9p�H|��3���="e��<����������� Yظcʷ����Y]_
���P R��Z���~���-_��qi=ڥ�\<1�j�w5m�ӏDѾ'亽[g9��������mP٘ѳγR�~@d��H�G=t�H�p����+?��t+� ��@Q�T���=��Nٽ"�'�����Ս���#��]'��)hG�>����<�oY�s'KF���9�Ѱ�%�v7=�:B�����#����\�vn��g��Q>ނiV�Z�<��drSQ��O+=H�KU��[O}�H��6������2/�| �ռA�C<'x+�����{w������WORFϔ���'����d�ؗ��Ы��/ࡀdS�Q�3�̝�NO:�«�<��	����ܷe֞��#W�a�7h^��,4�.�>뒡i�J�ϗ���o:
��t���K+����?W����gg#/���30�ʎszID�ub~�����с$�GƋx��Tt�����}r�W��
�~�CW@wc�<A���a���]��RN�M��L�EA��a=X&K����~;�rm��_�:��DVr�&s]��0<0��EU�{H �ȏ����V�x�-�W)ֱV���H�z�'.��u�v��`�c|�r��i�dZ���"Ot2��'����g~��]
�ֲ�(7��hz����9��B�r�	d�S�O��	#N��cm�=S���5�hm^�3��n+�FD���Һ��=f�c
�ۤޮ��k�b�p<ım�m�g<3��>&S���/¶�K��Oqb���nf]Vx��tg6o��0�t)��]dr�R'dsW啉I��l���z0ֻE6�pDt� bo��O�s�j~���x�jx���v.g��MM��}����B��f���%06^����Q���7-E
D�����j�&C6��q��f���/3I/�P�u�v�b�bY:T�}2�dx:��C̀;�a������
�0�ɾ�|�[f(ʁ���-���tm�6ߴ�����͂E��t�4�������,�&z:�=X������	8FF���E�!�Z	��j�������A��&�VZ�:��9����>�~�����}"��b�#N��ϯ9%�`v��^T���[�t/e��͙���y�'=����r�^�IT��3y5��`�<u�LoBAI�K��Mm.�.H���7�:���ᦻ�K�}�����O6��+CA�2i$��2CV�%��8�W�.��ߤ�Μ�h%$,�}����t�1����RJDm�
wlp+�Y����0�h�v������F,���!̯c��@�{�αq�&�j�K�er���x��#�P�l~��=ti~�^�_���݉\����&�7���T(ɉ~)���:2�b��y�{4��)qȐ�����F�X�%�&_�8V��;�<:{�E|�U�6y���ұnLӯ�r7��q����XY^�Wp*��y���ه$Ht��(�QZ�c� �V�n������n�)8q(�"<��ރ�b��Z4H3��������S�u�(���K������Q��.SF�(�ѻ�HNl�{ĕ2�2-���߻��0���Vu�mშ�q=p��K�Ұ�ke�|�C�}q'��쀯��Cj:;���@$&z����ߴh0t�Dk3�����J���~?��!����%�nP��M�Z��?~4���¹/�aƮ�J�팇�?�[������$��B{I�nܪdͫ��2��9Z�F�ொ��V;��|}���=8ߩ�q�Y�#�*�M���ԗ��c�9�0I�-(X�'`nn������L(��<i��h���*��1���{�%�R<�pn�65������>�ګ���dÛo3(pzV�5�dk~Qw�*.@�2���.�"��<�"���p_��^NI*h�hl��4z��&D3��H,ϺF��V��uC�5w��k7`q #���\[��Yo>>���'>��~6��D �S�;$�V����.�͍��u��m��F�P�`;ל�Y�_�h�.-���%S�r�:}+ ����3����Z���wSl�(�gSzA�Aq�4Ph��ڿ�N}���ߥ�ti��I��q0��Ϗ(�o�u PΫT}e'�K��S�HSK�*��=����e�,CS�|������q��o����M�$���p�h5@����*VM8��Q'm������P�@O"ܕ@L��zu�{L)���r��6)�Z�m�i��
<�r���?. ����;��С���I�������y��>M�b6%{H��6Eus�b��P���OI�ړh�2�j�f��D��ʡ��T.P������y�p�	c�o�mWߌ�O7�!��p)��"�"*����';����a�$���L�'��� %��tz��T.p|l��aWmWiZ̚%����k%Oꀰc�2n-�6��-2󩼹C�#q�1��bmp��9��YF�V�����̉(�l[{�I��Ôp����Q�S����
���F�����//�5���*T{®8l.k (�L���Aj���]�X�+��.��@��)����Ai������N���_#w4J���e��.�l�(������B�2�����r����N|;��1��W���ӵ��M�XD\�,5�D�8���_�[���n�_�;2q7-��>��W���^SW�O��<�T_8�����N�h·�/xA�|��� ����z�^Y��}s����פ7�w�0al/r��ⶳ=O��?���F}\�Wwaz��^^���s�8�w	�l��8�^�����Mz�w��+%�l�t���� !���V�E�{�`Y�6,>�+���85�{u�\�uֿD/��K��i���q�G����1l�Ƚ�e���7��Z��Q�i�{uǖ�S�6�gh�*����yA�(M`/6�� �C�$ΤxF��5<$�	_������S�9��1��U��/�%�_���e�1�	�K�Sn�Ќ$]���O��.^�da�34��Pq$�o1�G[&�Itw����,��ج��\&��`E�r����a�����y(�Y+�;����d^�v��k�,U�(E���⚯i�W^$����~�;�YQe) K�;�
�� �־鏧D�WV��"4��*�H���z��_WEV�Nh��O�ā�,
��?�� ��0�*�ii!�o�8,$�z_�}�ZB7b�4�ѩ4n��Όg��&Q�(�v�������OV��A�Ⲭ:+�֪�;[�~��98��|PM��6��hg�E�[J��	�f�N�B���	i�*���<�aE�Z�XDњ��-�.0)�'ѩM���w���#�@>�1���̿�!��8�=�'�:���/x�_���n�e���#�'�N�:u�!?!\��lșV���_�T3G��E�he�¥t��7w�W�hXؑ��Q��Y���z�R�����TFh�@��|�w�c�)(.T}΀���>�K�:��-�E�qw��H������ 'Q'��w�Mt����zSN�"�@�_�58��!`*so�|����-ԟ\��A���a�gڦ��C�m�����R.k�rd?j17J�y3e�Jb���sY�,����O��A|B�."�S5�ur�$��p��H� �QLVWTY��h�8=ΞZ�Kxi[���"�4�,8�S|�$�T�)�>�(����@�uu�i3��\ݍx=Q{�Y��3��u������e��2Q��,^�}��03���Q]2yb�K�C*"�	��Qt|%H���~���1�ogS���5����?I��P{�t�d/�s����}�f����o�!ka|��T�r� (���Se��+�H㮂7�)���u}4�6ș�4����)�w��ꈹ�{�����f����(���d#fg���'�n�9�k�N�F�)�QL�Е��?�3XF<��/$�E�ǀ5�����ޗ�K���6���M�:�G��=�a�U��{�W�ȮaՓ�9UN_0�|T�ʌc�DZ�w-�*g^3.�3����W<M�,I§Vq�W�x����N���7a�Ba !�E����r?��
��*A�껀3���B؏	DS���?;3��m9Y�F��=)Ҹ���k�@Un�j&諏q�둒��m���&U�ⴄW�\M�,�P;�݈O9�J9P��#%�p1R]����N?����F\浴h��*�rFD�R^��m��Q��2���F������3cV�+Q���{m��t�O��}+�J�A�G���D���T���1�*[�|���L�i��m��@2v�z�~׻��rY�I����D6��wM	M3�hJI��coE>�����zml��z�R����\���%�!ћwb�Y��<��2�gz��$.kv'RƼ���!��{�DF	��!�^w&�	f�v�ۤ��o:��"�K�3�����k��ã�z:�_�bEi2�ˣ�rMySʎt���Z�WYaܡ�Ty1�+P����؆ֈ4��1��A�.Fb�`�]���t��t�8��>w&��h�F˛��� ֶL��L��i}��[�?i��Ok�q'�=4�Wޔl�mo�s
\V/#(C������O�l��!�R\�_�S"���KIQX�(@�����cR����E�K�����#�G�Z����ODN{6yJy�EQ�>�B)܋&RƂ�o{1�A�9�|ȅr �M �|���S	�0�����Ta*�jFխ��;�F:8n}��[�A����ZO	m���L�k��RGzF�w��u�Ǭde�ח�%��9"=e�yY����w�
��"�+`f~�C�j�uEI��E���@l��.p:�eÎQ��&����0��+v�T;л��!r/�"tRTk7��f0�Qe��?U��Zl�w��a@�HT̨���vWXS��O)~��Ǹ����Q@�S�q#�i��t��!���9��I���*�lv�?6��H��.^%�[p��HB���b��l�m��!kk�W�8��b�Ō�ƜުwG��і�$��j�$0�@^S��Ax��4�h�Q!ml4א}fQf�2��=>P�'�)��$�����䯚8��}I?壠�p��z�8mIm��^�%x��u#/\�q�ZD�*��mB5�Z�J��~��zO.n3���� >�޺)�m�O(������#iJ���lJ� ��<��:'��u��2�x�z��V�X?
�R���Ƿ�YãtX�7Z������I�v�C��}+��;P����PS�4�R��M}1��!1�z�oU����D�fCȑ"��GI���t�m�_ٮL �&��+a��g$?�8Ʌ͐�ʰ�Zc��$�sR���������d*C<�M�Ǖ9�g� �j:3�;�G݁�l�I���e�|�B�E{���,9�d�P�z�n]5�k@SQ�B��9z>�F�!�X�1a�K�Q
=�6���&����`��?���(�A����.�F�y���[H>�Ǣ �K���l��λe�fOh�g4�F�ӿ�C�bt��Lg�AC)P �R	op�#X�4gL,��VƢRYϳ��owQx���f*��^f��B�O�%��!D����/2�������#Jy^�pT�L��x��f�S3���N)P�2H�Ƃ~��2��Lg?x��$�U웢�7����w�j7	!���ֺ6��qS��7��<�A�,̲�+g0�j	�ō�ª��E�憐]�C(^�F���^������W��)�GNLd������Gvi��"YCP~l��bt���+M�8W`�'i`38a&���y��-j�Ld����&��� ;)��E�	Ś�l��Ut��܇��I�;Ȕ�h�?��	���7&���S�P���2���x搓�5��u\2��0�.��� 8�+o�$Mk�\f�"l��C^�{�Bs)�>��.�vur9Gpu�۪��D�
L�H��8蕔��ۗ���cS��s�1��� ����\16�Kt߼�+��WM����\�'J�����+�I�ɘ���	�ڮ.�������Z�	�-τ�0��zu��/��Ѯb�?xf/�+�WH�-v����T>M?l��䇵�U?e���<���k�����3:x�p�
���wk'|o��Z�A�]p!�'�{�V��qwA��S���=�\��?T�B�~��i���v�����G+�p�}:G��F�Ӣ��[�W3�wn2 �1Lf ZVE�R5CP ��E�vcߜ=�e�A����#�W���pC�Շ�<y��M3� �'(��R�!�⩱�	O,x���.��0�
,�]��0��{2��c��-�9�� F�GU�L�K�la�_��P`����psfKM���ed���&���`t)p86��(t|�N�Qxo�-Ve�$O�-��A�&IV�u��?�z��r��N�kÃq>"�H���e�w����n9����3-cBϟ� 9�*����&z��A+jSE�T	䚠�ȼ�F\bߧ���dc�k.����@sv�-� �
� [
���m����m�7�S+��^3ۺ,�8s�Fܺ`��5�u��q�aɓ�
z�5w鼣#H>�w|8=���m�)�t�$|@��t	~2<^��C���S�)����=z}�4��mN��dZ�
y���-258	G³:	��C�R�{�V�ng�c#fcl�I�kw�8R��	�":)w[�ڼ5C���D�7Y*�e�F^	'X��l��gc�?�.��W��X���9�΢j=˅em�F�)�e�K�VK�ϊ:�t�
WQ�/��ыg6<����6��t���7^t���*���ݴl�.嫷���x�Q^� <Lo7�}���(�g��V%�ܳ��@�-�+�^2���ι�q8��u�1xA�npEST��ַs�*��ѹ��#�k�ͱ�\ީ��Af5��{�X�y��m]�T�τ	XE�ӬY�ì�=���r&A�"�j��MX����g���F�T���/�u��O�Ы�*sI���`̑q���\�=Y˦����!E�:�������W��}M%��)A���^|Y7�.)��gBXc��װ��I��H�,�����j0�0���PK���}���p���$r��B�UJM筷��6� B���9�`��8�$���2�+����	&�Y���C),ic�(�n�8���@;�x�k�$={!�잵���J�x?w�P���@�"��
un�w��u˫8��مQڐ�>i9q�ʃl��3"��Ap��	/���r�HʥcF�e�j��3r�톥��������2�����[>j��kS�@/��̾�P���
�P f[��WZ]j��l1a�]�z��hB�/�����yzO�H��l�s�t@ �|���b]mg+_�� o�j���W��= ���[:<��Z�5g�'�E� b&/	�]M��ǆ�P�tW���
��jC�P��H�t�AN��.K�Sf쥶�6JiK~��k��(�����8�p�f�K�rQ�,Pf���خD{�#�.wx֗�#ط���
*9S5]���P_�	?����;[�56�Nۨ'�*F�S�����͛���G�SV�.5 ��&c��7w���R/t�Z�Z�{S��������_���>'���K��!�����<a7b��ɬH�_,�v^��2�Zk�����yr�����C��rœ��H=$7��ڰϜ�1�P=U������\���K�TU�;pB�t޵�m?�~o�ra/]n�iG���`��02\�i/�O�3=C"�Z��&�mf#֔��"�.V�Ȋ�u;��V)!����@W"#���/�+�����o�ƫ�;RH�Wy��_[<�e%�3C���Ó���4vsL��y;�t�T�÷�����m{�<�ɧ�U1�lGc�]đ�0��U�Q�������cajM'����K
�x`7�Ǎ"���}��ޔV*:_Fe��q��ǅ�����������%��T&G����8�*�Q8�a"| V�2�ș���D�6�0T��=�����'e̹�`���)a[u����D`n�<�R�� ����^�_������z#֙�J�4�xxn�K>�7i���1H����� ��Mr�U���*Չ���De�cGT�� ;�x[M����H1�st�Zbx�}�P��4(���}ȌB��[&E9�n�d��m;{��6�N,e:�s���=�m02�<ug�4XK��F<3��M��"�ڌ8%�����~�J��z���Z�#F��X�TΚ�H��a���gĄ6�?,n�~7��%$���>s�-ciYM�$~��S*a.-�H++�1�f2y�z^S��|�͠Ǳ�D@�֕�fON�f{��[p���:Qo��鮲���lg�_��_�V㧷F,�F*1����=�z���tI�1G#Ԃ��Z_�3��K�i� �l�3JPU���K�|��l ��9p�� 3����mHKW����jn?�Z��Y��9�b�c͹�Z+
�F�i&}��'��M\&�� 4��CF]��0�W;���p�I���B�v46�/J�Q~kڀˆ+a���ܺY�D��
�`��E��N���4�3��e=���+h�)��2m����=W��}��q����B&-�����)�b��8�	�l��5���Ɲ��):�c��NV�9� ͬ7JE��붯Ⱦ�	v��u =�#���*#��d�Xg=�>J�!�F�6��BS�����w�l�ګ�v��=F�Y���(z ���Y�T��%��K�۝]����]�BI<��f�y�g��8��L@�-��S��D���Rа���mӓE�񴥃�!c{X*U]�M ��w��O� ��X:r5p]X\�D��j}�2��E0�v遮�RX��I��~�\~�{��l^�N,����m��Y�z�Ơt��.���Ќ�.-$ͯ��a6����O���bOb�:��ͅ[4� %	����f+A#��n��`miRG��&B"،miZ%�����E�y�?V�a��-�Q&�k`>
�s�&U�[,���������.�mc$�_�.�P�^֔�|9MV��M,[%�=��0S�_%���ir ���;�ź���S�m�3 yf(�t3wY�W�^KB��� Q�B��Dܓ.��E��������y��T����F1��tB�`/�8�<J��	��/�4��?�a��
��.���-IfD�O�sqN��i�����R�c��>�gw��P��<�M��x�m����*�D*4���0㩨��A`q B�̠m;��ެ�b�Y��	�����|���j^YI�G��~1S tc q�m˹%��Gm�j[���S�7�or}�ʙ��D���ÚtGR�8Y��ڗv*�I��o[9G�Ae���8myy-[�fXK,>���yAvg4����L��k:9��S���<i�x!�(�"C ����v���c���@�We� �Ｐ�/?��<����yR/Ĵ�[��+>"́SȠ���D��L �vx��]��x�7�ri�dOFE������n
�R����58XpkW�c5�!��jҡu[ww��|�,�� 4��Q�gϙ�S(m�/�,�S80�}��3�x�n!�,��Ոx�ΰ����*�Jn6��4h��y�(c����\��+W^�����Z�Uь'M�c׆ꋑ�AA-B��|����Je��V�U�DZ��xߒ�w��5y�N �Y��Z���Ǖ��vB�`�;O!�ߋpOF^�^s�����MzV�K��8����Hz�<YHa�� ju0ɗ�ܻ /��#�P�1��b͛�_�l'�-D�b��I�KH�*��V߶�H���@���vaS��9�U�+�LaM�\Z�U�Y<���v��o�\LƏ[@8}!�#�T:!-�O.l�{[��J�s�
}�3Tہ�*��\���O ���xis��
�����QD43, h�8��$T��h��a0� Ä��!@W0�ɳ�c��0:M�󔁑Ը�QC�i&���;��]��8gB�uU�����.�v��z���ڻ�=�	�(R-�K�&ӭ����N�,`l�(��WߖF5�n~dS_�� ��k������?s��xE��.v��^��֞!��T����:�9�Z��cr.�N�C�-
��G���^�[�~�;aW�
�zp>xs���^Ht���%���_���k��@��K3D䔫ӯ����fNg��IW�.r��C�.��v˜�ߤ�51�ɞՔ�'ǭ؞�O��@7{��X�1S��MJ�U�H���^)ʂx�%�2�øK>蒎�;D	,��Tb�n��5pV���p$��DIV�v�wE?��ҫQ	���[����=��D�5Ŀ9,ff��"��Jr��^��_�!/WՒ�|�wb��1��Q��I����,�N-�gݑ��JƔ���+g�[sy��~�����R���K���=T���k.���iuU�[2ʏ�tQ%�[� W�n�il����eǿ�/�6sl,`���n��GU
`�^i�合��T�U����$e0�Ƹ��u�7~�QF���6jOU�~C^����ڌ|���pPD�����k�e
+Ԛ��|G��+����J��ݔ���.U�K^�=B�S(�yϓ|Ӷr�h3�SP@X"����9��L��I��V�� afȻ�sDIL���y��k}�;�����̉DF�=����T{)�^�<�Aև���NG���WE~?�i���' ĀUR���J%&Ue�Ԗ#��������xW��p��xEAW83�]��U�bs���C���In^��<&�0ä�O�Nf�Xt�ϥ�����ݨA��-W�:0_��k�
)�Q�2�%�N|]|�iS-��F_��i�Jj��,6R[�l���B�n����+���t��:c���'���1k�Z�K04U �{	��t�N!4¾���2�dD���.|����`#0l�����	������NJ� ��=)��#	f&��j����S-��'��)�a'yk�)؅�IP��ؔ_�(2�m�M��	��&�[�K~yd/�b�ϻ*�1m�r�U*��C>?I�%�V$� 6
�Z�Zv���=��@���/�ï��$��-n;�jPcx[� h��Jy��.K�[mvY0,gK�M��%�_�o�~�Z�u�P��n�/C��fV��,;�r��H��e~5����He�vp��-?� �Sr�I�P��]�ǡ��hu�|�,�g�g���{?n�fW�d̤�.�x`(����\7Q�m�JB�`C��*�5��He�2؟�݊Qa5 �f.Y,[�8�*\�Y�i��� �VI��=]���),�>o��a�:�-����d��j5H�h��@��K�ڹ\�ץ���k�$qhd�BqPP~��w��?�-��V�8�C�' ��^D�� �]�������8�c�K��2�����H�~v�=�U�佮�;:�x�L�q��/�P�+j�f��D����0TxKޮ�7}�N��u��Z��9�յE� T��.̥KxEhQжq��^�����`6���e�O�����dS0�m�W?�F:1l4#卼�|���|�U���Y��"�tA$�D��	F���u�$ه�V�0f֓�C��ME}�`1�L�"������)?^@X
QT��C3�@��78r�����Ƙ�Zۋ}`��9f�lkQ���z;�(��꽐�"܂JƯ^`����`1]�6�u*4SH��h�	*�YD8�d���=���i5��"2w�R?<r�=ԶS������<��w�K8V�����=��p"܅*����o!$�ArQ��zKF�d���v��q�iPP���VͬL���°���K��)(^�!��]�xD��I�0�QJ��r���c��9�1v�e�;��G�R�7_�3��'}Lq8��e�U�%����J=�R
P��|�,�O�uʺ�or)����<=�YS�������Q�	 ߺ��Y8#�Ajx��cQ�Q|�f���������w�<Ԛ)7Ѩ�p���7���pI�[5���j!n�wpQ�� :�zUuE����=�;�_XdW�Y���1����p�U�~tP�"�c���E;�>.��H�J�MO�h�c@�Őo���;{;X��h�<d��A���-VwsN�:�s�,�U��c!P�}������/y8������%"ws��q�]����ȿ��b.��a��rx]�:����.����H��rA��/(:6�bJ9E:o�W�~��BP�XQ�?�x���j���Z?C���SR�7�S����V̎*��:�a�܈N���$�ٮ貑O0�eE���W5��.ܘY�[H��6�4��f�N,U����+�ձ��x.L<"��x���"6��%&�b+k�-�!E�ܔJsL�L��Z;}<�Aty=0��:٘P y�Eɞ��2z�k1�t���Ւ����>r�P���0(�>&ۭҗx������W���D_p�9���}��K?�v�#�^Ck��D�RT/}�����`�Ⱥ�9Mk���n�K��6I��������NL�96���;�-8�r�A�Q�a�"�^ʪ�#���G_~�ZE@�y��n�ט����e�����r�ZI��<������ZG��m���P�"Y�k׉yଶ`ۙ���"z5ĆIŬ��i�� ��Ї�j�le4�I�&��:�*��A4���zrKGm(����������h�.肽���N5|h�;h��:����1-!���[=��[b*ή��G�]/�O��2V���̌�J�>5�ѽ�*��~ݐq'��j�g]�x��Zֻ����w+##�+����b��y����ԧ�#l�E�X���-5F��Q�/�LT�y���J![�H�w�l�	��ANKW��������n
Kj�>x³	�T�%��SB�e�X�QI[�xX��a#jg��3]1%V$C�#x�g��FjT���i�_��A`1�U�3�p�59�G˲��f�*���_�O�7D�˄v5$�$���hu����t�CtH������ޠ������7���8Nw|���ߧms{���Tn)o���#����C�fK3�R��SP�ֱ� ��������u��ҬP0
;�� $�%�di鴣��H�s_H��Zs�G��G�_���ڄ�@%D}{ �Rz �?6��`���0�{��^� q��D��o����?����7��!���$cC���l���"��
r=�J�j���L�s�N���3TD��e���7��3�Dqw��U���Q!!��P�d�	$��Y��"��V7t�u�{�v!8l��<K���O�:�o|��k�+��2"�����T���xXo�6��v�����]H���m��ٖ3�e��Q�ۨ�_>�!��������Ns��7KZ�ֆs0eOAS&��~u���τQ5t'Ș~��g^ю��!���낵	u�s����w���sﴔB$�g�
�f��q����]��e�9�;�\�Ndw�+�z���6�ȇ��p�3��LS���+9 s_>�˷��m���#�y�"w'�sF���37�҆z���:@͈>�	Z��	�� O�j-n���:W��`��n�,c�;�� -#�զ ����?L��̌8�����4-��|��Z��h�O6�'�4���S��V�!���-���g�so����>ҭ2&��Ce�1(�"a�w9H!�l�|I�]q��Ɠč�7'4�9��"�LHwŭZIYQ~��W�G�eUv*��;3(��#�,������0Mb؅����E�7M�B(`�|�������M[Z�G�u@!�k*p��M���|�
����V襐��������G��H9j0u�x�2�O\^��5f�s����i37�k����F��E���6�QC�R-E�)�W�SI����!��KLK���]7����s��oBERQE�ٻ+����DL���ִ�۰�����=�9�G>F/���ՙ�L6�������]���V1pz�fS�(�WE2�h\���՜�7L&�{BP��ڍ�� ��]��rYb*�-!FX�E^��t>�7[cz����f�^�������.��>�s���|J ��ȴ�
�hkX$��F��[0��l�+��}��&H��o	���v�l+���h��̼�(�yg��T�VO{�iן�K�f9�x�%�pۋ�?�|
�-��k��_7IzJQ��Ї��K`��K�r�uĆ��D�$[��3Ж�\/�O�T��p5�i����OO]�Y��"���?�9�To=dp��iL�"���"}7�:�gr��>���� ���i/�ǋ]�S$YN5 �I|o s@�摂��è8��QHo7�2VHD
@�]���P��Ru��fn��)�^NeKS�\��)�ڇ��̨�q�Y*�=фox����\���rwn[kj@B�*wh�5�0��E!i#<���:�<��9F���[��E���:$
%�\4ę��U��5�+��q�M �E<h��dL(�O����'@�d��DM���<ڱ<|�*�E�x5�oyWx��g2��c|���́W��\~mq��S_>�'Tc��R�x\�M��ܶQe�%�%�� ߧ4�K��v��#�Wd��m{�
v<���BU�FT&''�5<����3ٌd��z5DH@˱�N�jܣA�"��[X�=��
��u�D �{kz��޵p��E�8j�=�?��r)�.#Ӷ�@�h�t�ryoE�������]�J��T�B>����
5� �y|�T��񉥺�⫣)N/����%��X�}ut͞��+�'?+�C<
�>��8]ao#�fu5$��y��+�4���%E֩C��W�s�m[UE~��F����G� nE����ȘE&k�'�r> N7%[n�v�~�v�erN�dO��_!\�����!_�$� �_�'դ��\FO�4ws	����f�v�tH�vaq�7/l�[�9�y�C������v�5�!�k��1�^K�,]C�����f�@b�Q2�����'��Bӗ��%(��k�Vw'Q�}�9`�<Y(nKl�ڗ�q��C�j��ĵiLw�4�c �C� ����ƛ�ź9
�M^�n��®�<p9�����hc��v�!��6�7bA��זJ*������$�T���P:�%�#����K)��xmۇ	L�����~�Ӻ�^8c���IH�+2J��x�R_҅��a܉�T��qIk:�!���R�Q��7��l ��T��W~+�(k����M?4�D10�·)��97�Gpٌ��t�
_�h��N��썒[�t��T���'�m~��
�v�-\�,l	��@t<Um�g}�+ڮpnpm�D�)	�~m�?�9=p�/��ȶ���b��_��ِ��W������=�7�71l/i�9~C�Gެ���*~���C���گ:P��2���_�T(��o�5=+�ԃ��#
z���,!�"xK'����%��?� �2]6g�
k�5���Է֝K��8���m���6����"ReYh��8�A.
�tv]g���ن�Ͳ"xFz?/L���iB7������V�ĨY_�y&p���\��@-��I.e��(����=�<c���!���FTS��G�2�D@ҝ���Oy��ՠѶN�K��+�xs#c��$5H�\	�� ������5�^v;�'�,Y!*�(�&��]��������� mەC�k(?�P}np�1kJ���'$F�u�t*<���Kq,��L�~�tՕNsy�����p^ ��hg�q>�<ͭ`��z��T�һ����5(|a���vA|�j6g�F(@�K����g@|�
�k/�������a��!R/$�f�s[yX�ЊPI����V� xA>�T'�N�^�0P^�U�Z��H�:ؤ:���#�-a�R�@�>���*��{�kF�C� ��%V?3m�k�A `�Z�5 >��Y� Դ냕7��C,�%.�E�:\T2�%a����}�w�܁f-<���=�c;-�~��q���P�v�Y%���^Fw���3�Gv��{zg��M̓�uZ��D��rg�"�����R���U��#	��B<t�0?c}���/��k'�զ�:���pqv���ְ�z�F�����e���璷1���Iվ���i���k��X1$̮�2�湧�Lk[�@�����g��.k�Q�� 0���^��X����զXDu������e�Q����o*@wsS{��Ge��H�'#nEV��SŇ�&~*)�b�N��c�6CG�k�=�`}�Θ��bvp��*�{�<���U�"��O�f�3(%���{�1!0U���vϟ[���}p�q�@�d�/xv'����Y����� \���ҋ�����Y��CvY*R����:�~& �	&Ct=R�B�]_�'b�;M�� �]���5�4T�����{ʷ��nK9�N��n?�|�hg�*���_�����@Y#͉���/#��[�]|{&c��=;W��-��&��bO�ldU	�KD��&KF�^���T=�|�����a�-��jÕ��J�!X���۪e~��l3������V�'6�/-����?����}�b����R�~Ɔ�Z�	#�:��<B}0�TH��Ò DHm��.Wk��Z��>/.��� �N����.A���)�!��W�E�xq�2���L��J6=
���������L���P�RPU�O���<����%)�7����k�6iiͥ�vϟS�ߐoG��hri=; �J0wWKV@���yJc�ީ����=���@�M�6��p.2!d�,r|S�ɥp˝L��GV�E����I~�Z��<([���D�) ;.F�$8�<C3�s1���@���1��3PUʢt�yA�/Y��mC��*�7ܢs���s6��mښ�❟$�FB��K���Rʤ�OK�M՗ �q��~F���l�$ ��8�K����fV�zo̸�q]�	�o޻��[�	b0G��y���.q�h˽>`O�0�
�b%W��5��T�����]1ۿ�`��=�Xq;C{3t�Y���׎A0	��oA,^bC�*൉��O'��F�~�P����X��l�)�V�${[�-! '�V��k�J�(SL)<w��y��4�E��L3�a	��u#n�%���K#�!t5]�����u�%�X�YLf��^n��O�(�(^g���)e0��iG��e�&����3���sȳ ������$W*s*���Z
A�v�U�:0�ǹ�Hn���сo�W��'���b9�X�,��I�#��cܴS:�fk��ء��Sx(�����������մ̮��ʒп�5����$Nݷ	D��zR�B�٦a�����@�H�:t[~G�fZ���c�5|�|�O:�/q��#�P^�ʸ������n���@�St W��g��h���߾�(Idev��`b�tf�ǵ���eJ�0Ʀ�a���O����%a5چ-`��;7z?U\`mFO#Ƭg�����'�U�T(�b�e������� Y��L���qO��|��C�WL��,�'��܂S	����-b�fNO:U'x�?}� ����F��jE��,;������w^���_����W����d$el~��Q���L��ަ�1�q3���S͖��\֔�!���<ޛ(v� 2�퉓&]x��Dx#N��V���=&S��i>���/��#�p��khNWO�+$��]qz�Vji�h�f"#
�Mک�-b	�Q��ʍI�߶���x�-��Wղ������K ���w�^Q^��U7|'�-C��瀚'#�p��F��ԇZ�9OR�jme$C��4�Qz��Z8~�E��R����1x�P,�퇀�,�ȑ���o2+5Q��$�3g�6��f�5���~*w�R3Zݩ�\��G��c{�E�%�1�@-E��Dj1��bx߈�/\��qĨ�'�"�+��-��/`^ҡ8)I	LsɀDm^g���hL6� �`j�����NTj�Y�9#�~_��Io�(��z�햠�ɸi�O���}��8>'�N��!��N�+a�w*�(���V���xs?VolV��/�kŵ�F�v��	|cN�W��"�F�˷�>�A�՚P!��T���C������g�6F5����f4��>m"�����
���QC�?�������\h��G}ls�u�/�N`W��f��z5�Bu�s��@.�@��G]w^�K��������N�5���G�D$��W;���Pΐe�����4g�s���uV��6�
��i�h�'�$�=k�#Ӛ�I�z2��W�ɂ͢B����{��5�PK�ԫI?�@��8���|n�"�S�����^v½�����A�x%���C�w����I��I�S�Ы�Sr�%�F<Fma�f��ry��ո�������*�y��s.�?�?B}+ �+��2ԻRE�%<_���MA�	�;Oi���<�"|pD��l�z�M�B�	��U�tPT`S��k�Dxs�~�����X���e�����uw��x#Cs��V��?�Y\2Lё�%��4��	��s}�����E�o�#����M�07Gn2h T�ģ�g0�#��'ޝ�7 :� ���8�MR�ܦ��{��)D�G������^Hj|��ĲmQnCy�%�f��+I̽V���c���b%���}�mg�9����?�y�G��s�1¸J�;3n��"��C\y��l������Q@�ޭ��_��֯u���X+�tU*����:�6��]K<rB�F��;2�u���,[��Qb��p���r��{)i���{��
��g��Au}	�h$M���Ts*ا���t�r+iw��&=N����P��g���g�w�Σ-�ĥ�e&��ş���ۛ�%��~p'�23&t�6�1�d��8k�ڭNZ ���/��#�5AD���w���A�!��hF"Rln5x��/�GI\��$W��ry�e�ߴz�B
��&��v+���w�FHf�>�-����D���Ւ�n6�4��w݃#P�+�`��tF8*1%wC�wz84��K~i�ꪖ��I9t��x�g1���d#7ٓ�t���]���T7�߁���A6�W�k:!)���w�醾<�v�X�&�K�P��h� d����7�T�i�*v"�jU.�#�5������C_e��P�5�/�L��ey�<EǍ��$��**u��D5���˹�53X��C�����BѸ6h�6��ءgʿ���ኖm��a���/;����#ަٶ���s����P!2���! �~h�^b4Ѳ�J�s?E���6�S=SX,�A`�JW��T��[��π�����S�m�G�U����&�f��-�����L����|ݳ�c�a�q
��T��C�0f�>��=P�'��<��es��d����\�������h�F}S� �:�$+�k�7�]Jd������?��1JA#jE���Ϳ��5
���33b{��G�F��h�g�cw�R����z�y����G�i���b�Ceb�e�+W�U�M�.Z�r�(�Y�Z�nX����J ����td�qQ�U��B��4A�La����l�͜\�[���P�fs{���ǽ�6� �m��#h���OΙ$o�sw(�
~ru�I���=���H���eaM�;���6Vձ.�߫����$"/f։�rݘc�\��Α�y�x�@-��L;{m�|BpQ���W�7��.g����0�Z(e7�D��O�c����{����**VAz�Ϛ�:��Y"ɬ������cʚ�)E�z����x0s�'����hAt8�E�J@8���F�`E�b�~�o��bf��6��8>3�����7��=o�)y�?�c�0󿴵�1�#����Y�o�6�&>Fhޘ4<�^J� :Kz��?
�AX:�E���SpBt8z-�ytJ�}�=����8��f
74-�*.������T����aR	o�H��Ke�R�O
��U�5�	G�d�T�C� ȇ��7,ΠC_���T*�
ø1�4ɘ��i�؇�w��o݉��<�nX��a?�S�} �+B�T�'K����阯/�dpīR��{��GZ@	UV�{��C7rEbhrTF�2�<�h*A��� j����&Z
��\;�F��L(�l��v-)��K�V� �ߩcb����QF�'[R�5��f�=��g'�!��mb�@�;�-C_��NV&�A/Q���Uoy���RdwvA4qB���g�ah�P�~��<�*�����W-|��Q΍���e=g*��|K;7a������z[�d)Oز1�]�Xפ+j��?F��	T�e�s�3�pچF�4��w)Y��]S�@M봀�m�(j��b+�ND��?��?$A�,� E��ϢZ�6	q��?3(N�`�]U�XH> e�h�s�5�,3p�\��Sϵ&�ڴ9���ç(3�v�u}�G�3�@�B�ʍS4W�P�d^r=G_�L������v���R��� Ƌg���mFGM�΀f��ň{>��`ljr!���C�yM�M]W��>�P�7α�޸�6�� KT}���z��f���3m�n���ɼ!�=OX7�8�F���ـ���TA.��N1*�6���A~|O�ǧ��r�l�XcJ�d#q&ЭLyc=
�	���F��+>���|X��E��N����fm\�<QJ i0�*��1��M܂/�`��r�W�!�Drs��=�	�������®b��!�pC��
ݨ1���[��4��$�"i�.�����p�7k��L�)����_a�2���f��e���#G����.f�b_Q�B#�9�R;~��>ʲ�s�!�qM�朞�ڶ�����)�J�R�rʂq�A-k(�j����R�t6�,o����y �~��+C�2�Ȕ[����l�k�m��gyW�t�.����� aCW���������Hb�xFF�y��c[eC�}&ݞ�))0΋��a�f�/7ވn�&��:̱]�|Q���BK|�i�8~����;��t�C* e��	��E8�柼�g"Dw��������tP,�UF����Q؅���Q��%$q�� �Q��NǩX�(�^��%^�H���Tw_�@�ΫqQ�w�A:9G��M�>z�.X�A�e�r9���>zⅲ͢�p��R�/n��X���\�e�.�(z�p����4 Nǰ�a,�`�īy!rҐWV�L2#������z��2Gy����-�<w�����6�ByP��(+�c'����.#�.4iϯer���;h��������*�(�g7��`�!���rdǒS� �8sDu�\<=Q�r����/	���\�4HB渪	���Hfj}������΅%�^�5�zLO��T�p��	�r�)�?Cw��4�:����đS�D��0I+�v���& ����5]�����;W�:(�P:C�kl�z�{�
>,z���I�}@�-+�T�q���������pR4��!Jַ4Τ���S����u�+a�d]'��F��/a�D)�|qEu����ް��`������i�Đy������)�����4͛uR��*K&�*E�$[(au�}�k�V�d��-x��>*q� ���X�(�V�A�h��� ����]Vr����#�6E��ƚ~u���s$[���.�zM>��v-�z�@���d�B�#e%�n�s�8��r����"B��:�-��R�M٭��Vg��̛�F6�8�a�u��}��������z?�z]�����R�}K {_�0<����3�nx#3ꈓn%:��ݮ"x%{ꁦ4σ���I����vl���,��rg���/��q�\��}+;8�vk�����_�E�F���׸&<�[���#~�%���p�d��'�M���%�.s��)���j������B�y��`~����DTMI��'�ĺ����ヘ��)	�&�vT���(C}�'ղ�kL�]s�
�Y;V��ӐZ����L7h�dz{�P�t-�z 
���lJ�V��t��]3&-����꾪���"�+���b��	89�G��E�х�I��5�n��@t��g"���Ď���1v�d��G�]m�H"�.jrH�ӭY��	�@���P�,F��_������2�tCEΕ5H_+��B	��
�) �j��1�)ӐAe���x�H�йfm���y���t�W��F�-���x�]��ª�a���v�Q��Ź�:A6%%8�_��f_���>)�N��
6�݆h���J���5
���G�kn�n��Wr��ݼP�=�2�9Zq�t���:���K��N�@�x�� ���u��e����9����1:�-ps���DE�mA����`āf[[�T
ՃӪ�l�Bcw��
������[�9���
���S7W}����xQk!��R��Q`^�]d�Iq}6O��L\-��]p���\v���!/ �b��:c&�������ҩ�s���>��ۑK��K?{J!ea��ΚRMw�Q��FR�DD��pq�1�$� �<@�k/Z�F���K��5�"�><�dK�Y�6`�V&3����?<��8G���3lت�LB�A�h�����`�����D�I(Ƴso�yn��^n�mju��C��Ե}B�A���A���c���DZ��X_����d�P����8�����mz���tN����e�)*��,A^D{����<�q�CI��� ��f�l)�z�aJ�C����2��e�z��	�̋]X-p��Y!@�~�?w�8yjմ�N�^�{�쉱qH�p2�xi�\t����U�ԁ�ME���<��)2�N��>�{��c���r�\�z��ܡ��C5�wZ�l�V4ހgߞ)��V�q�7�'���������7�_C�§��vז\s�fo^H�8Ț��*�U�P��dfwr�U5ezSSp�����^�*7�v%�̞t[����&����&�cK�~0{J���%��&�Y�4�AŌ�1�[���<���T\�}I�BJ��Y;�N������f�!�Ӿ ��q�D~!�nf�|j����o\���&���HԼ����٤8[�7�k��0�e3����8&K���[�p�I����6B&��g`�ɰTir%2�l\E�|���������DE�I@����k�uop�+��\�ӟ9�PH��~�ğ*1zLq"�AS�_u�^��J���^�͖�����I��@��p�~����a�q����HH�����-K�͌�L�Y����+n��+���\�,WZ[���86X�Sk;���i/�ٽI���S���S���(��w�$�Hu�Vm�ϤX���6���?�~�C\�l5���Z����B�R�Ի��<8�V6��$�"6�@¥'Rs���+ؽ"�b���q$
EN��q���?~#�l�oo,�P��3���`Q�b#�(��7gHr���SE��(x[@�۷-��~<��׸�0&%m�}����P>v��9�!AN:�wW"�]����?�(��`�NW�s��Rb���O�ݎD���hV`���z���
�H,�>�ܘJ�@�{Rq)
�X-�֗���2�������dY�UU�`E���H�)"�"���g�;r0�����8�r��hIR=�if��U�%BMv�w�Wy��wV�@'J@���Y��!Ym@�r}��K�̪�D�8hc�4���V��A��\��r���#qa��W�����Aء��Ԑ���t�$4�=�t���á��D2y,Q�����;�>�R�|x�m��DF��]=HRb��L��|m�X���z�n�%���~_��빫�n�R��9��O�񵦣"���f��x5��p�u�m�-��q��m4�6�8��'�.�_Q2WA{�a֑W��k7�(}6�졮�����x�y�#+��_t�?\+�]�2�}�H�7�b�qV���:��#�h�����$��mu���E�^4M�c
dVچzw(�m�tJŏ|D�FaD�v�]U���F�^#b�8u�rFf����发�~����4�oRr|t�[�č,�q^$�omz�e�i�o�$�\%�p"(
cm��!(MO�u��8�����oa�vؔ�4gIj��j���^T��b��<��E�7X*IN�H^��3>�(\ﴭ�S��g�5P�B|j!҃�J;j2���>��FT��,��^p���XH�W���#��I3��Ͱ9�+��/����P=��a��X���p���`=겮�N�l���ֲ�<e�̛r#��q�=��(�Yƍ���,ݲn�e9�QU�QɦW�lq��ӏ�JA��uk B��1�dP���+�ݔ�1)z�_��Q��;��B��c[ip����8��P�$v�"ک�ӹr���6����'5�(u��J��+c֣L�)�3c�#a[����rR~����G�y��a�6Bl���R�X�������y`25���T��������G����k�dy��4�`��Ԑ�G��3�/�$C߳��L޸������9����R��d��gE��!����B�X�	��{�-�@k>&���j/�h/�BrZ%�uc����N�2�a��/�+�k�7ޢ�OѾ�=>s�ݮ�B}<����:��2W�2D����p��i���Tw!E�	:J��N��KhS"�ɠn#�J��Pf�}��pJ��(��U�tT��飽ΠCyC
�2��aR+n�b�i�KhBQ�ؽ"ۡ��*7x����*V�^(�Kz�-��HH��?���DPT#tX]F��w������3�6�1�b(��WS�S&V콛*EO!�J��<ka�8�Ը,L��'D[�w�)I]_q�^2��q[_mφ�0�Č��h&��C�����ai�o25���[��P���멗N�N�ʘ��_�*�c�qE�wb\���N�Yd�q���(b��Z2�k~�R���杒}	�^㊪���'>��,?�?�R�OR#��;o�Y��<#-Q��D������%�F�
�r�`ϩ}?d���,ѫ>�R*����87*NJU����Gm���Y����'�|9��.�^�qIA�7D�K�g��Ɯ�]�߂xߦI$�1h�:��]��Y-��}Mڇs��_�Y��Jr��C<9_���\̟n��n����Ґ�ɯ��e�>٩� 4
�]�a�@f��L��ʟ��q0�$=g6dj�:�xOC��g��Q���+�/�d��#�t!��PI�M(��mhb~��MסL4�,YZ����n�a����ۻ_�Ϸ#���J��ά����oAx�rNָ���78��¦� ���!)t,(�n�&��D�Jݪe���CX���v�������ց
�U�q�S��'�[������!�Yh��Uy�� �f�-я8Q�4t���#�bX^w�`���6�뭁��<�J��wy:��)�x��ĻL�>�ŌD=�3��i?g?eQi�ʢ?p�@#���5$F��ԟ�MY�f^�����M�nd�%@X�鏾\Õ@rF�g>�-�K�DG�V&�}��[��s���9^J8�>���z�P�v�M��� G|���p2\p2����a�-��c1:�*�{"m��E��n��0JHf	=lh���\콙d��{���Г��]���9(=��
��?J!_�%�(�$�����hŔᬢ�KJ���k%|D>�̅9g_h�"C��LKwm(�c����@��Q�Z��<���}�k�S�P�o[E9@j(����.�!�:,��l���%
㼈SZ�k7�6��,jY3O��CME��#^��:6����;p�@f���R�c�2N@v*���ZY_���o�z��w�M��g�S[���֌/�ƫ/�(+����	Z��ߢ8c�~y���B�qPD�}2ë�Y�m���k��}-���Y>H��h+�Ń=ڲ���A��>�-7vyN��q� ���xe<q���4��4�G�y;��tI����<ֺ�Vc�CRˮJщ��<��K=V�	�Uc��T)PM/!ł�U�ACZn��:�*.�Jr�F%v�W8
d�2 �V�}�Y&�l�l���1xjf`���Xi�Cԟ����Ƅ��ҽ�`�uH��X(df�O� �E���A��9�v�}!�R�T��"]c*h2�i�4����VmE����s��0�7�خf[��[UE��bcZ������.3�2�A��Q5t�śEI��/�?E��XÑ�ܱ7Z�z���b/�LWqXBT� DYWy�^+�+_HT��*���/^GI��Q�eiء��2�G�ݿy ߦ���g�3�}ܾ��w[�*�����=F�	X1�fTM����f$� uk{p��^z	��z��W�d~�J��<�G�Q J���5d��շT-��H�:�=���/ ���JXR8��p�&Eh�̮���u�j?SQ�_������<�Hz��#(W���Q�=n��L��s}��4�AO�sG �a�%y*��.ʙL�:�v#:���1��6�2��.�W�z������Oc����^v a� 9� ���N�=`�\��:h(��7���g(�~��g�03�����;vy�L��%�!)� �A�eDޱ׶P�{�8�s��d� �mK����A\��� �����lښi��Fc� MІ�����w?�p����[)L�e=�U��7hbW<��>��C��I
�>��F؀�Z	�]��US>���-C+5������ձ��.��(a�M~N���0"C�li�o�U��Q�u�C|S�K�u�K4���c�Y�wg��tV6yui7���Er|[�.�7�U?jf��6���ѱ��Y4;�`�����ly���f]fD/�E�=�rڅ(�l�t<���E�N|O
��;��:���LL�:`�k@�벁߫z���A��"��-� ���r���%u��y�$h|��� V�ђ�u'`ݗ1.�Σ�ܛn(�9����gl|!M�C�ӟ��� ;�jﺋ���n����!�c�O�	MQ�2J�Rj��f�R}������ʣ~Q,(�,��d�����7[%ȺX�r�Qif<3�j]Դ�^A�&~���>���Ԇ���X�q%OG�*f#��J{�^�d�T疏Y�U?�!�Ho�k�w����OȽ�+����6&I��\�|=��3�ŒR�7�Cg)��5����F��­�+K�v)pj;�2jJ�#q��.P!����a�T��Jx�X��ݱam>� �����œ��ki���̌x���Y�r�����s��D0�l����yY�l1+_�A��6�ynL���A���,��:r3||Ty�]D�/�!�j�N�xz�Q���}�q�yA���"O�����Dn���Dji#�D .�}��%��̡�bxȮ�[���N)���94M����<D��X��p�Q�ЮYx��r��+�L��j���qZ��Y{�|jk���W�ڡ&u�Jx� B�^O"��Q}���>�#f��Ƚm�����7���:��$��Ί�+<�	�l���J/J��UT�����9��)��esW�E�U�,O�)4Q��κ���nQ�����r�?ع����m3�V��"��pkV���z6!� �h��wK��n���o���߁6�����"CvtG �%i.<��yLdB�LՍ��Nx���!����d�K��įS����,7�p���������b*m���U���'�R��oZ�۞z8�{_x���8��V�A�<�ⅾz&�g9]<�����m껇�U�k�l����77���m��a��匿:D��d��fA#��X��]��=#����.�G�a������(���/�U��?�&�Ff�X!��_�4E�$�+}���y�� 5����立��(5xh��_�cص��E���d��:�|��k��$�埝G��`L��{��Nk���S@��L�Mv��� Ո����n6�cV�{[�qE��(��r%eͣ��a�3�	`� ���U>�G�I�����Щ��'��^ifބr��Go��GLi��@ONkh9;��WS�G����F�y�o�N��1��\ΊUύ���e�U(����C0I�"��ɛ��h�	c"��}��RK��LĈ������޻"<4���Q{C%��K�*މ�ţ����2c�{������/�: >L��}�(f���X��1x��'�i'��D��鵁P�s���7��f46㔚�:,�r��^9����~����!v)�خxF_�41���m� �51
�z,�����LU2ϑ��C����wv�y�G|\Z?pE�S���5����n�y���}e|Ss[9q�f ���4�<@a)@�s�rn9��xZj��\"h�N]�N�]<r����PZ?S"6��ZߕOeg�J/�i;����� �-�	P.A�gq^�5IWOzN�Cp�}�{���l�b�o�E/c�# ���.h�(������������ ���;�rH�8��:�~n�@�1|�H����^��������U/�S}~:�:��cͻ�X��!��:F7�jFA6˸���-EeT(�`2Jqް�@ gh��Z�;�kǦ�ˉ��Sv&���J�_�>�á�%DN��ql
�>>�ve��-��c4�gABXdo����T���]|F; qjC�Wi~˨�Ob� ��=��}����ȁ ��uy�����,Yl�Iy��Y���8d�'��Z��J�}����ϙiN��>�߻����`*,��9��.�N�^��t�j��ǡ���m�$�{�@�Er���Y[�	[ic���{p_�<d�@Ne��6+k�����i@oB=Ʊ.�Yy!-,�tF��^��[L�����.���`���7c/�}���� �k+	����"i<���-,���U~=jV�2|���R魶ꀴ�o�asS[w��=�$�ƬY�Z�p��4Y�J	;���wkԨ�����$����G�1=F��H:΄�8
�!zOza����{�"+��f�=*� u&q &a���%�R���SP��V|��@�S�E�,���xeu"�/�W*�oqG�����vQ���}J	�EL�m[V!�lٙ^��}[�kķ՞�Ru�ls,Jm���'��Z1�^�|��~�e>$��Z��rK�s�W��ֳ<���?<T�+�5�s�5����zeQs����9���$�&�b�ME�;I��t�t΋,�[@t>0'\�a-��ٓᬏk>c��V���w1N�<��0���i-�^jZ*�+@�A�z5��7�׋�{{�s<b�G���?f3�e&QgRJ�j�Hء���@~�O�
���H�'g�`w�����m����&W*2a�G�r���&�x��'��.��p"o�(a�;
6�&I3�2�>��J��p��W��t{��}z�\
F� q'����Y����y�j�lإG�
	4�'|~�����2rJ&��LN�:F�`<����[�4[�NdO��j͠�V��|�	�y���4��a���<(�Ѣ}=o�`-�m̏k� �<��K��G��cLS����JE�Z���kƂ�\�МLa%�c��Q�w%9��#.������h�B��1��H%�l+���mJ[��������M,3˶��e����������-٧��G�v�$�'$,¾���a���"�q8����#����N����|��v:�J^(�bm�_��*y}t{@�B�_mѓ�c.�XH �{s��ԙ`}Ŀ��]����>�Dqt0L���*ͱ���Ab.�6 �W��KJ.��Ux|���3�����V���F�������彆�S�;��1�{NL�Y�$�W�Ӹq�v��Ʋ��48�Ȑ�˭�?�w�=E�(�bN)A�w}����ϯ�8��ɽok��LF��ٞ���@?�y�������:u�ѝ�x5�69�m7���D�
3�( ���a\��^���ۓ`��OS.�ov�$'jct��ш�<dy}E�wߡ�l�6�Í�����DI�e�Ш�EZF�)���n�*I3�P�)��Xf�pB���bvJ���)0�QhP���k�1��ft�.�Q�}��Ư���$qN"B�\)�;��l�����-��:
�'
~���Ԣ)����@*� ����0�0�c��=��dE\�h�e�Œ>/���MgQ&@0uT�g�x_�y�-�#�y&�{ਙ�fC�4e/<e���o�U�(������	:����K��郑��e0�v�Q���f�w�1d��̡lW��b{�C��9#AHi��U�m��T_LB7j�

)���d�h��� �}P6viA���o���n��i�_�1ޚAYp��+}�0����'Q߶�/Ď\�,\J��Sٲ�aP��IzBD�>�������&�d|�c�X2G4�Z����������O�� ��L�,:z�찕��X��D�@�ηb<����;g�@1���0���/�� U�'C?G�+ѲM2�t��Uw�����׌1K4!H�� /��Xۨ�#5�]�~�aJ�U�J>~3�#�n�A�#�W�mm�J�j܎,�gw� |��yE�^��X�X� ����7ri��ءiÜت1��#4��۟���;ٴq��}�߀�z�iR�ks&��R	�#	(���K.�Z��pL����X�z}�W�:�wH�æ����&�@��h�\��4.�ӥ�8�������j��zi���:���L��;��K��Q�hp����n���v7�+��%���9��8S�������<@���M���\j��!��<��@"qce������t-�sD�	2Y��s��t�`@0�|U�^=� ��y�����w���V�V�4+�³�Ǔ|lH�s���+�@3:�6~�I�e�����z̚����������-,�0zA� �u3���*/3�J&���Y��r`\!�M�Ep�2H=$���Ȣ�8%�E�4dw��
��3���z(���o#�糺*4�����}?�%G�cq��7�l�����E�d��[��*�n�(;i*��,�7"� �p���a-,ٻp��F��a���j>X�X�)R��U��HH�����d*��eP����6��=}<�#�U)��ކg�1������E
�k�Oo]z,��Ȧ�m�V��f��HN����%�֏��V���0ǣ�W���T���K!n)�	�%�����X��⢷7�*$,�3j����gI�X9��Зi	�O#5(�S���>�j��t(Ed:��%"�^��������H�|S�h\İ,�۞��<v���v��O��q��gw��@&i�a�؞;0q���p
��X�>��bP��� �)� �Ї5x��9�d�r�FD\o��$I]��Cm�@�뻺N�J��3����X�-�L�m��,ƌ������aKn=L�q5=��gi_�s�EqZg1�2T�Y���N:e��Cg�{�R����SޚR-���z�Ɠ܄��L�������x��P���T��Apq6	|z������-��v̀񎫦��X%���%x�#]	��8��s�b=����}(�ˬv\�=��Y1�0	��O����$��\n�CF����U����m����ubۃ9�r����<����T���[jp��<�,��K|�J�՜X7~�E�J�����"�=�פw�|ß"���R;�
��s�	^��ǂ���T�������^�>�}�¬`��z)��~��E��7UZH�Fa��V~�c�1�~b�j_.3@�ws�~�:vZ�Ҫ,3�#�Mx�!]�V�ޑ1�{�ڤ�^p��DG�-�0��E=Y*h�k}u9z���i ��r�<�n�W�4�t$��?P��[���+du�qa%��EeZ�m�Ab�S��������Q��'���Ɂ�z�Sm�o����\�y��==��s�ËT���ĊJf��BP�r�
J(D����ְOL�����L`̜)���+n��u�U�Utޭ,*7��B���Bc,�q�*�
����:��I�GIG"M�et��vd�N�|2���D���#@$]�(��c�� �0���
ј�O�q$�B�O_[=m���u��8ZL2�^��	k�)a,L����}�s�y�=������n|��z�#�g�Fn �]���P߬C�I	�)@L��G�9�_�)Tt?��T���"�tǂ���}��`D���ɽ�.qK�cO���y&�x4n����n	0��,S��� �p��'����x�+��촻�v�-�
��y}`�1�-p��U9�(P�_5c�"������]��y�Z�1E���E=��K=�m�Q�ПUXJ�Fΰ(�� C(PM<-�߂�D�f*Ha,��ۧ�6�����"���]�Qi�k� sи����Q�z/u`k�=Z��;yrk�H<|�9��vQ�A"�8�C��U�4
m��W��z��ĉ�ޟxL�ܹ=r`ڮr$b$�]1t�ϑ�ЀT24�W�kb���Ie�ʐLT�&�4_0c� �f�E���M�>���mB/߬�V|���7�q���;Ш���X��[|��^h�j�K���=��,��f�Z�bч��ԟ,��(	�y�3�xW�j�"�}x�tI���؁��ԋ��$��=��.B�/.�Ax	.���%��e���!��qBu�9�I��h*� ���5�����r�� 1��
 x�<���u����)�}-]��Ys΀s�{��OkC����!E:$:�b7j���wV,�NZG�(i���Z����E�;�ʣ�E{t<G �4U /�&���*6���W[�>�\l�o�{��g-Y�[1r��Y�s����u?ue�ÄOo�"��O@h�!��� ��R.�Qg��9��7��s�ien�e��3,ʽ�S��4U1�����<�f-ߟ6�fݽ܇�VA��@_�����/�8�d��J5ݛC5�l�_�V��Xǁ���\76�.�(�����d7���r�߄��S6���r}��hX�μS^��kQI���"A�`�J%T�0y.yE����cM��cE3�j.�����O����wG�"��؍=T$��X�p��+F �n�o{VKx�P��q�З~��
�� ����=P�����f-~�bS�× �f���K��{g��ݶ|qM
j�*K�#M
�h_�OJ��C�`���0�\�$"�Q��P��Ҧ���MD#j�H�	�"�锡�-AW����oFV�#ʶ��U���>v��ǲ&���s�V�ߣ�_�kF�$���<h��ۂ����Zi�t^��s|.^��c������)j��0�
�
��|�ژ������S��E�0���K/�����=҈U�d5��YE�_��?0�}�qM��y���.��iW�e�������?1F���e��^�eI�-���~�>��/Zi���� $��GO�'z� �?�Y�Aoc��1�Upl���R����}Y��eT˻�4
zC�Be�_(�7��Ӭ�����;�v�isr%�uj�A)'݂�)h��X2�[1���p.R�Rb���y�NW��>���3i�B�>���&y����<�$e���9�f{T����Wd�vo�]*i�R�.6w�r.w����%�����a�z?�3sỹ�A}5!
���Y�c.P3��&S�I���cl�$��]葂U������kvVܙ!!���ʰ��o�}���8k�9��t#S�ㆽ1
u�/�����Jo��	q�N>���в4M"�b}7 w�"4Fbj��*Q�m�|�xlN ��$d�'���n���bg�?8ހƽR�_c*f-o�2��ڽ�.�\�;�¦-IW���2P���
�E
h�oЩ��j�9E���1R�g���a����00^�����!=�?xZ���W���I3�����c��٩��oo�	^hB>�\X��K����*ke�6�`]���j�&�I킓:���C���lA����ܷ�6;  �1�H ����t�G� �*F�I���8����(c�<��G�&��:L����[��`�z]+Cꦘ9��P��M�V���%�@��h�ߕE�$��{u������墾�'��5#���`mu��i6��z�!1	��7���'	�"���dk�h����xJ+��fı�N�����ݩ�._�#�+�3�|a�ȗ=񦭪{�b�+�V�����a:���a��rϠ�R������ ��0�%��
�-��\�i��-�S�s��u��K˖��l�cG�<ղ
�����U��k1A	IS*7�S[�mF�?�\�;J�~��a���s��j�y`��s�� ��rF�e��d\�K�{����!�ݚȲ�!z�D�i�gZ`cO6@�^��I�8�p/yxӑ��}�FbL�<Ϡ�qF����ۅT���׃�2�2�u�1�N;����4�N������F�����T�|i���[n�沿�� ����-h�����q�|{lޮ�]e.o�&$;�?x����&���I�f�������Iþ��'���o%Rl���b�\g��RTcd/b�a�0�*�8�l�cØ�e+��umef�{�Å���D��~~t�Y6jGL���c��gz�l[{�����L_�\+%En�:ݽ���,d���^x�6�g@D�����+'zGr_T���oM�i3@��+�����X��6H��a˝�{����e�*_����>��]��b���W��<W`�} }J.L�q�m#a(
E����z\z۟��wJg�P���Y�5��d �{i=�w���k�es�u"���)}zV1����ִ��K���2/�T�b)�2l��	'���T����M�H[����,~:V�R�)G\[���z�?��
�5}0+���V�/���h</T1����LȺ+���^X���-Vu����>��e�����Ua^-s��@��D������=��sp�|7EF�|d��3�3p'�nHR��aCB�ܔ�Y>���A�5�k�VJ`�dr��[�Φ������9q~ɸ��_1'J�p�κ�{nR(��Q�UK��$~n������4�������'���l�-��P"�a�i�.*j��1]2�%;?!���M�5�(Bo�p�S�4��sc=Ww�ǲ���3����ab�Wpہ����l���1/�O��2{{h����.�[��$�q�G�a�ޞf�KT)�9b��<p�m�b��i �����ys���nٜ}�1����H��Y�dHV���j]��>.�6,l���[T���{�+{`Ö�D�p�m)3��.H~!�ǧ��S1ᖥ -�ޣeN�/��V�<�>��L!�Q�+s�0�:�p�2m��bwqc�������M���/nZ�aCa��չ���l�I�\ �f0)a����G8��I�z�m&��d�@���|�e��	'{�#kh��OF���C������-7����R�3d�4|T������5PS���1��5�0�^?��r�&��G���ٲ�؇�Ri<#h��<��)l�����O�a>Ʋ�M��s8DƢ����D2��'�­��Ղ�|.G}S�n���p%�y�n6S����KZO�>���	��qrU�_>���%�)@W��G� ���n�� 4nH���0A�U�6i��O�CfY��^M��"V�%�t�M�pH8���g�L^����C�E;o/�ڂ�PX�-B�6^k��L����`Cm�x�7ñ�9�B(�[��<j �@ҘD�);��Iq܇lw��m��i�pж�ǵ�$���O��
H��R\�J�ؙ���NC��;��J� [p�CA�����ń8� 2B�1�4�6H,�M}>�1Z-��_>:�.B [l��)�ـG�/
{=:�K�^VS�vr�W�ЯEQc�#�v��4`uk�j����'�@�Cvj\)(N��i��q�y�ing�MsP3Krfε���f=)H2�{�3MPC��J�g� �ޖ�r`?n��۹!X�Wp��l���<E��r�����]�l��e��l��H�*��9��SJ=@0n<rI��0�����T/44�����]����O��#_�����%�M(7���&�wH0�8����/iB�!H)�p��a>���J��|9([Jȶh�e>�����@`Np*:�n ˛�@��K�0�����<��XI�t��5P;P�,e�Wq
��x�#۶ƨ��g��(����r�~R�z�{e�Pө5 n���#�������զᝲ�7�ǈF]]��>W���͚�VR��٩�~����[o���*jT����7�m�h�p���:�*�xC6LEl���S;˅��V�;�����ʁu���R9dq�"u�+����}T���r@x�V~��d�#�hD�s��&>�2���(
�Sfv�G�ܬU�U6�9^�c�� ξ{����ꊍ�:��kt4�����Ĩ�]*ը �h��5,ܳ)���J�oݕ�D�(�N���c������a��0�[k0߽b?��m�����r�֦�vd��8�x�H���E}�jC{��;�F@�y�6�V0ژ%��k)�䯼��������i�N�mC��*;��|�%C1mx�����"��0���rX�[bqo����m�Y�fmc��D�HM�8*�R'Ĝ]��tol�e�R��IH���"��o��\�ֲ���'��S�:��}U{���W�+-�� �q(�3�_�A���r� ��뙼�B��4��@:4da1� ��+Q�ˁ]���O��"Q=�=�yE�֏�cLW�!L5 &~d��C���ea�ٿ��_�I�kˉj�����:g�չ CcA\���h��ߑ9��8�J��,5�S�`��$�����%���1�����?�o�&��X����(f�W�3���ۓ^��"��L���
��.��c���1�dH^�d�ڦ1����i#�z=G�	0�e�Ku$pQ�i��o�k8��V�@�yF�%�����A+Ql���2|B��V�i���?�e�<(�1qi��`�{��)�K$��վC�||
����vQm�?�ȒH�S���֋^8��0�5�}�S�RW��P��4���bJ��ErM����m*|��SPbJ1�D��@EP���#�-��O��OL:��L�&��PJ�q�dEKOVF�\�'��M�'��$\�`@&<H��r^�,�[�s��6E�,��J.)L��x��PK�q�RU����;hi���Z�蠊##���;�g���:to��� ��G��u��v�݆�\�`���R
p��������WX�ӧS,U<�ҭ�h���UU�K*`,��L���l����S�j\��~�ĕ��d:r����	�[�A>�TK;U�*�	�6�5��\�8Qąe���w�]�F%�R�͝A7�x�V��W������=�$D1�&!�5ݑ��S#�2�r�hF4P��U��,�?�$�+�)�7�c����7a��9���y��{+q�C6�k
̮c������,.ӭS�ӳ?C�c��ȟ��	�#��eǌ�����0�n�}�E_ d��!a^�R�S]#H���?k3�GM�#�D�F���b�2Q�kN�V e��O���w�a0ň���I��Ro[7����ݽ)z�n/(��T�d=iZF)�Ȩg�"�j�7 -���a)=��3��|�����KP
�T}���
�?�j4k�p ��<��-�W%���ܲ�Zi�b/W���P����U�l$Î��P�H��@vR�@v�j���O�eK�Dq�{��3g
4��&綇nzt�O�}%S�������na��i,�)U��dϠȾX��F�lߊ�D"^��z��WƸ�?�%WntSG�D9�Y�)CUh:$�O�`$�� ����)�����F�T�&\O<pE'��I6��?8�b1�EN�X��O+�uY��]m7�n���xkpX��wg��y�Al՜�0��S���a�l$�ph������Է&,���`˫�Oag3�ѫK��qW�L��e�y�T��@5�%|���"~�_�3�Ě/Ih	$\D:"���Fy�+&�jN�2������11�/���Q��#)�9�А���ا�t��H`�R��K��	�������w�4I�HxNN���+χ$Hm�)&ɇ�H`�*������ѤF�ȅ�'������Pq+P�)4��K� ��?�6�%	Mф�v�F�C�ݜ(!^�8��Lu|	�ϒA@1u��^ S��6-oە�y;LJ�c���[y���{�Y]D =&!���F�>�S�����PK�%���*1F����gr�p�ܨB�ߍdO�R��z�Q�!'�e��� �iU$��� r�V^�X{�,��A[��8������ʹ`�H���F/,��բR�u����M�PC~vG���+���w��ySV�8������SB_�?�z��qҙ�u�U�	����uE!n�j����Zy1������k*���0�:��[�x!�˵~K[�8��CЖvNZ}��3�\��;[�1?�D^O��E3Y.G5 �4���:�Y�K��VE�]�=�6��9��o�|���ٙ��*N��YWW[B��z��f�W����i���Vf�A���OO xyl/��=|%�'�H��ʝ�fKh�G?a���7�E�1i)�c��\��T�:�.h��.�tc�63pN`!򡖚V�Oń�-al��8��O�ʋ�wu�\����9�P���>�D��]ߒ��Iė:8���M�Wu����Ҿ{����+@��6��a�j���#pEi||\�v;����W�L���ګA��).�ú��COɖ���mî��)H����!���=8�ۊp��U��ms9�ʫ���~�j�^ޔS�c��v�l@����h��"�s�?I�J�<�����~�E�A$��|'.B�����3�@!>�J����5 B-`̊{4�z����O��%��b��M�~�S�����^`�g�+{��;AQj�\��)%އ�{zS��V�5���Y'��v?�N�tV��g�����=�$7(��gi>�_8�T~���y]�%�=~�O����&)�&gG~��-g���#]��]��R[%ϩ+^*Q>�?҆��$�2���� _��a�Ҿ��[ 0!�'B��O���l�+�>s2l�����3=eO��6�m���͗͆0����%z�#��-+��#�~z�nl��i3�w��ƃF2�sWdA��-P
�U�%����9�b����D��s��i��M�*m��!�d!���.�N�#� ���a�y�,��U��o\&�[�{��K��{��a��6��,���5A���π�b�2{���=ɮ�?}V�R�><Y�.
绫�����I��I�oM����)S;�tm�nm��y4�����?�)&Zِe�c�$���y�b�;o�0�?-��а��
���ɏ�a�g`�j��ml��@�<	ۋ/m#������e|)*�گwaN}�����J��<���p5
CZ�I�H��i^���:�KXķ�7�� �m=v[���?]����e%����U���r�����'�%R�}�k�-��͎A���lO�U;v���"�����*�*�����2�<�ye�yQ�����1<�cq�N��RS-@�O�
�{���3���u���:��B�0�6s�f�F��y머5�aa7Nx���^��Y���;/[P��V)�5��F�P�*2�yq�gh��z��G{�`��Y�4�X�5�����T�Q�Q�׏���v�[>� ��3�N2eJ�$���Ů��SG�R�t��i��/�����Q�Y Qގs��Sy��b��Zo#]��y�l�wut�Ν�RocY�R@*A����z-))���:����o��<E��VF�䡣�AR��F��ѳ�i��CF��l�.x�s�F�ώ�ekQG����,�����71�vcq|a���~�H��i�C��a87Q�Ftǝ�T�U��&�rr]���;G�3�����j�3Mg�'�{�n�5\Zı[0_�1S�ۯO=_��aB� �%`*�ԘIA$���!������h��2T�.~�����og�M> ��赝;��
��O8��gPŜ�+ٶϮ��F��]��ܗ������	�F�87���~ vМ F��v�Bы�7<:չ�j�8�'���i�z�Ȯ���4V�'�S��|r��g)9];�1��c�K?{��[F�Z2�S�`$�Vy?wf8�ơK& �������E� �.���[�����	�ݥBi:T��z܌��eV2�n�lwQd?��R�A�=똰�+dd�i	�dKQ�9�ܰ\8�H����9Ƿ@&a�y��R�t>n���O�@P�c�!|�L|F�tT��W+vB B���l%�lW:�F�[k86d��&E(1�pS�+�R�a�(]��ɒa�L0�ʱ
no��J��� �ʫ��Ԩ�C�@��:%��Z�e���]�Goȃ�z$լ��u{�W�~����;���s�F�ZHq&.D��� ~~�YN�M?�����ij�F����J���x�!��>�,��T���?Y^X�� ⱅ�?����>7(�!L�Dbn�=^��H���" lb��t[�L"� H��t�h�rT����j5a�e�F�!��6/��m&^Xp�к#���?8���d
���y�S_PEM�bf#��,0�2Χov��ŕQ�ZT��bb�A��?9�3���i�o�����	<9;?��?�f̻d&��y�::��<[�vP�s�I���ɷ�/�Ic^��T8���Ѹ���Pnվ���������G�ЙI�;zϣ��
۹S��u��@� ��w*�R�{`J�*��1z:yeOo]��1 ���~.���[o����'8H��y"�qͿq��p�<��
xcQ��F��f;ȳ�f+6��xya�*�: �Y�X�_��O�	+j�Kw�z��{���g��(`�H�V)����F��`yY�a�%�l��qK)Fm�)��2��4z.����J<&�� �|a*�O����0JĚ��Iݘ-�ߠކ�6�����+��`9�"m��f7��W�c|Òn��;�+R��Din�5L�h���`�YS-3�r/�)/�W�z�K��0�=�&觌;����@����X�WTj�8 wUF2�VT�s���'��Ǌ?H���n9�iL¬�YN@`� �3� f�v�v�W	���_�)K�J�P����C���H3�fЋ�+<�9E�C��K��'��BsX�"�:_����a' �n8x�	���H�N\R��E9�2bJɴ|��7�Y�k|�)���`���=�h�9�[T@���"����O��ʰM=�_lӱU�+����=Y�t��ߍ�<,Q�◬������2��*o� ��O��'��Z�6x��AC����(��]�z����1�#�M!)# �Lc�tA�~E��023��;�S�����O4�6��?(��Æ�uP��t.��i�%ː���|À����)����L6y��9�9���o �����bi��T����A�c��{���v�.lg/�ئc�헣�;�B8 �&�L�ĀC�m������@�π�����=�[Ք�<�r�����䖣h��4o
�C�d4�0%`���������*��rd�B�6H�Hl�g�r�F&�o��U�@�̂e�o�G�H�I�q���s=cȆh0�EX��ϖJ�UBP,��u�K�B	aң�g�n����ӭ>��a��Y�!���A�N�S�a�l�̴?qzH��h��}i.ܗ�+�>D���rx[�
	�ŎT`����L��W6�����1�H���� ),�npD_��<�7{���3B9���٧��o�j�_*����'i}rUt�|r�Z�1�|4M��S98r�蓁<#����s+f��b̑4<mr�|zH6�G޷�����"(-�"�k��j�fF���¨�a����~I��h�P]��/s41S���9�������k��X=�i^j?g5��� '��'��TD��{�H�Fרw](�,�_�Ek�����P82�m�4���t��OG;�b��\
���u�c1�\�e�|aϋ��� ƒv?h�O-:oi @��{�.N��a�i����U-c\>���m�%�$P|�~�'�q����Ms��!|S�p�~t��/�l�q��� B�����)�%<�� ������g	Lp��m�9���<����F�ۉ�Ѻ�-c ���"^KD��D����C�O�%��OY:�]�2��!�5O6�<�}\�ӥ�,*4� �k�k7p�,�$�զ���N��.�֞d�2r���c&M�'�D!XRY�(��v���g���-�W�v���#쮥�w%�ᓿV�g0��p�G�	�Ǝisc�PԖz5�q���2%}�y`��M��M��f��̈e��K_�<gR!��~4�TNF�G�l�XR�o�@"����`����y��ԍ��~V��B�>���h�/p[4(H�I�0��/���/�q�DU!���t�=�!���,�\ky�E%�*�껑Y�xx��q�8����p33�,��	`0�f��h���Kx\MҨ�h$�GY�� ���KyR�{lS��w�qm���	�'��.+;5�]�F�q�kau��ؐ���5W�C�_?�|���⟱'����q�84�hO ���}���k�����գ�~�C��𜉇�j�5�TkC�No>u��j�M���J@(OY�`�KwbN���(��)���v��#]i6��F�6�?ezx��G����&J��gQ�\}���P���P���I!����� ��#��l7������̍Y���;H��Y��L	��׫r(��� �������f�ދ����������Ŋ;�ٔ#��I�SI��e����:ѱY�3Ƥ$��{��Y9^#�m|;{��~��Wd��{Խ�,#]��2|8]CW����7.c�Ó�LDhs��Ӆ~�Df�D��X����{�cG�����imj�C�8�T4��I�$.8>2k}���|����룡.έd4F�$3�'�i�n(���%ߥZ�q���c���8��Z�J*T����Σi�j���tb�OwA�{���S6�X�;EGakŉeHB`���O�zR+Q	����Nlҷog�@�7�z�9�pD_V*Af�x�̃fK���W|�&�Ym��e�U���7^��X�l1�&�p8|��W�D-��� 8aN�����Kq�4��T�RMt�x�e�C���!���
���Iz;���x�.��*��V'��D+�$�cx|p�
YΛH͉Af�����)&���%��J30h*h�uxu��N�30�.� ,���U���}��hV`��C(��h��$i�����o#�Rm-��ʀL-�T��"�CK��ȧ��R��81C��iѢ��,���;��ݱ��f�V�	Y�%X�e�3�������,D�y$N�W."J��駺��/Ē�������]Z:�k.h��2H?W��ʭa�(��i��<��?�G����C�g8LhZ1�1De����+i������%��%������F�6e#w��`�m0ah���m�{r����Ks'�@�&�~"ί��H/�+q����0u&�)3��E����5�3�ivu2��v�ܤ߬(q�
=�,AѴ%�S�"/���gH�,��%�p����.�>��i�Y_n����o���#�r�N��[9���x/�So����D7N�b�G@�����8r�d"�K,�O� ����F�*i'Ӟq�To�L}{�&�T�	Ԡ���A&r�w⩅,�ܛP�\O��yn�T�UH��]�q�V|��ѧkb-k��\���̜����}���7���#���p1��瞕������.�������φl���Z�I%�8 7���'�G�)��gqu�=���ܿ��l�s{N0��	���7B�N�3i����y|�D* *�
�5,��r���t��o�ϐ�dZ�4�p0���!�4����/�q(;S4�{	�q���<�ڮ�+XQta��j�g!X_3Ax��K�6Y���.�	�%1%\�����Vi�e]ȳ�'e�"+����u��\gY�鏛$[g`v��$rs��dF���jnɧ����^�JmL�ν��r��^i[�HNO_H�-�a�����X��r�h6�5ճMw���{gUq��%�h�P1e%r6��iM��OV��ZU����"�Y]��M���-(YD6�e��e=�LŅSZ�ć�1'g���;��̌f۩ݟR�j��}���[��jR�+��J?5ga�׉�V�#~�����<D�ʙ�����edW���Y�4F&�xrepT���Zt��vb0z���l��`ZU� c�e6�5i"�/-7����@�nm��,�?�e�Ӗg���9���6t �L�Gux�~0	נ�/��E��x���`�Y��	�u�xBv\;n���`�pU��}�x���t�
j�#�۳��/0\���pk�.okt)�����Y}�%q����9xEn�LO�?�U �tEW|P@���-!~#?.�U�۲��s(�� ��!|���Dl�bk�y�� �Oa:m/���&��-�d���2�/Je�R�ڃ���p��,�x�;"��W&X�sΞ�, -�,������5 �f��]й�M,�/���-s����A�!�8�#`W�<�E;AnL�V�iv�d?͢����OO֫�OM�=<8>l��tܒ�1�l�kwA�7��M�=�)C��d��!�B�~}�f��6D@�_��ih>{�r�8B����rx]
��L�����f�!�{ɉG�Zy�~�p3�1gϹ��|;����'�&�OU�])@�^��G��ě%��4�TS^��#�M%��?��AX_n�G�f�9�|�����0��W7�Y����vh���tMs=G�ڌ�RUf��2n�ę�-�@kS��>��bYfd�Sa9�t��[�;r^mQ�r�u��.��G ������ܿ�/�Ē'��*���ƶ���^�,A�чTۆk>�IH�����xiAA4+A�l�Y�k�Y}�C+Wa�(SuI�e��)��;��P2bl21s���Q�c��V#�G3�.f[V�/�a'��K��Mbm���i8�'�T:Fܒ2��ZӮ�������^������r$��\@��1�s���������V��t�f�R6�"<�g�h��[4�U5^��A�$7*�KIer�JSz��;j[N�>j����%��*��^��Q���D���S�v8E��)&ԓ����_�\֑�,�e��Q��@2��W����}"|7+ޣ�_%���3K��Ǆ~���4}�ƍ+�%�c��$�M�#i���0�6$lA�c������^ ڮ��4̧�»��ߚQ���!�)���f#F�*d�}dL�=@��	j5�/J�wtS�	�Y-��D)ퟫؼ� .�?#��P?�4��eB:�u��SIw�ӶF<B�o��ǂ�<��տǨwi�h�D��Fc���x*_�؆�M�R]'j�oP�z$bWB�;�v�������z��nK|���Ύʹ��_�yQ��vؚ�2���D��>Za>2�%�#�����'z_��%EYx�@T��+lf�Zhj؁MAz�qχH-��e�!���M�;��r>����EB� �}&�k��q���5�3rf���a5�H��=�z|`�@')�(d[��4J_S��C�lo�+�埑��Հy$%u���*��،��~jVР�3�p��	�˗���	���E#b�D����w����A�ҧ|�P�D���>9��ċ�A�s��3��P�	��: ��j���ύ�r�ܠ��B�DP\��6���yw�6�:QWE*Oe�,�[�͢�=��[�T�v��fXk
ҝ���Mʻ6"�;�n�
0
<C���<�{�zV��ݬ�O�ԩ�|�����Yy�:�p�d�	��3�P�r(��ci�HR���f�������	��B�Q,� �(�ĭl[����`j &޲%C�4@խ��O?fh�)�����;Ѻ~�U�U:���{��������@����M'�Yv�	:��Ca]���X��D�����#��9*�[�~C��dZ��\y�Q����|
6��T�TI?.�F�c�{�I�� � �������Q��=���a�����RHV�Q�bu�ՎHQ��g�TM�B1j��|�Z������v�]zw�hX �q`�"?l��cx���5x���xH��	#�QKN��y�*�8�l0?G����aP��,L�-S���FP�zE�P�`�KG��TAfn�����"8]N~"B8?7�qJ�K� %4��b'�c_�I��0�>�fhD��#��P�`�-NȔ F#�qn����@�!k�p|�	���4?1[�|H~bO�1�6�36�F�	�w��
Wu!<�����Ƿ��<h1Nԃ� /��U-�
��pJ����S^�F�J��gRם��2���{�|S��OkW,�h��7<��L�f�w�p�*ee��_��^��2�r�����qF[3K��6������JWu�����&�ң*ȓ+�]�j�AP2@[�c;%M��2l��o�~���Cw| dp &ۃ�	��t#�:I��<�J0,�{�&S������7�ʔ�#�D����z�ۄf�V&�`̦P�<�E�]��xg��H�;YA� '��(ǭo&M�������s$�Nl��\�Ѫ�m�]	RN��i��ss[M�I�ߕP���w���3�K`�iΖES�*�k�^�7=��0DB8 T SQ��i����'[�"怨���8%+�Ҝ��g�+KQK�{�8zQ���u�D��h��+���
�� 3K�փ�����۸���<��6R�x�;�Y9���}��b���T�v��\�S,vʃ%���$f�D�� �D�0֬���?	�oe��Ϧ��Ş����ë3�t��}З�!�y� ��+�����k�����@R7�j;����W��T(�\f�S�r���E٬�ZWr?఍���z�
�L��is�1�j=I����@]�F� d/N_�Z��e'� �MH8髵��7J7�2�z�j�5���G_�d|@nu�hf�*�m�~h���J��,�p5�%�}R�px�5����
����g��R��L �-i`B" �*��/iG���S<�g�WJ��WI��!��+lu�[t�J�U�F�K�99'�;-9��6/�v��~���B�>~|6�V��'���z�Ui�'���S�3抳o^�eW
���A˦��f�,��u�HL3Mc_|�I�!�<�/�x��l����x.�Kzj��Ad�
��0�2�m�U!a��_�$ahS�'ѓR��赧��S���_û���\'�Sƃ=�nQ����a=������
hKV=�=XiuB��pi�ś��B7�����_�"�|�u9#�yמ�"0��M��������Bc�d�w��P����~e:Rm�ˬw�����em�a��Q���\$��>=�lA%�W�}y�b��<�ǖ��C�iln4/��O~��{���d�P&�rStB'����c1t�����W��ᓼ����u:�+�V�_]�ډ��ˋ�}7��ߋ�r�$YY����n�[u� �H�W��j�x�<�����;4݁f�;��J+S��ܘz�Aͭ�z�7�/{�3��W��/��MN�eiZ�|3[ѽ.fo1x����#,�N����}YA]�~J����!�;�����%A/>���x���K�D�͊0��7<ʷ�2��F��`N)̈��+��0�����d�+3�v�3x��Wȴ� ]UƘO>7`f�����fУ<�w
�Z�]������
q��7e�
O��\�1T��v��C 
)Xv#%�n����_��c�G�xI��3����eRa�,X���@�+����l]��'�m#�M��ҏ�#sH_p)b;a�{���� ʻ]����1H\�BswUL�nn�&���� 2]t`��!7RjoQ�6��i�)�kj�4��O:ꘋ�.Ω)��Nƾ�����lkR^Ĳ����)16��O���	q��H�5:�MT8���Y�9�Gq�΂����ה��iY'�eG��+/B���*U�ҳ���|EgV���!�y7���E��$���<)t-��C\��7��F�v���n_^ε�P�p�{��y�C/�4g `43_�H	��N�hm���VȖLh[k��V�3��l���k4
mH�R�"e�Y,|���ѹ0���$��c��*;t��ߕ�(����1t���!�gx5T�6C�v�w�aJ��@f��J\ʽ+�� դn	Ӣ'�����VۅVZ�'_!B2ρo�I�7a�er��Զ[36��$���q�e��B,��R��Th�&B4����e��v%����Y�u��-D'w�V��{ןI�+����2G|>q�&@�� FW�&h��1�&��e�a'p��!+ʟ�+�'��M���n�h"���rSp៝(P��R�f��x;���Ǔ �X�e͗�̨�vn����ԑ�%�4��3�[�i6�㯵��]��'<ύ��F�_ȓ�>D��nݽ�z�*7#��!W_���{�@L��A�G���c��~�Ń{�.] �`���$��[s�*I���ʤ_�,����#��(��,b�����S,��W�QѺc��u��l���C/��qÿ�i�3"�1�v�pfB�]����:��Y ��I��{6�|Lb�z����M��i�	/� cNGp�K�'1v�
����OG9�z!�����d��A;W�=XgFB%���ڿ�Q�+Kem�y�^���Y��li78�h�q�#)���S0��U�/ej�����D_�,��M�5uz�[��,Y�.��֠w�!5h�fe���S�_��1VR VB���xB9��v��9�{�����"���E��.;���E�����w5/Y4��g����N]��Yf��ʺ�����'�	e���eY2�=��*���[܋�g9��\��B����A�Z���N�`�`1�M��4u��nѺ��$�M��ް�G[X���4��3�����{>��5�$ۉ�� D�_~g�H��Q:��(���^��~e|��G�«�L��}V�#.8l��'rV�Ȳ�ȣr��� ���%2l�襾s(�y��#*�C`��j�T��ꡰB��%���JL8B�SN��ԛ9*n�"�AӼ��҉����;��oh�:QH'�鸋~e�e����o�Ƨy��K�@0M��r;�����KȑDy-��}I׉�7؅0���]}m!�*��� qZL� �ݗ=� ���*���Xk�~�H�E��6�}i_ �:*qHw��h�U���Hg�X(� &���(�=�M����mUO��3}��/����m6�7���"<�=mmdX���#�j�Tq�4�D⬕[#O�M�E�� w�s��0��`i�s�ƈ\?FG�Tyj�D���칆ŀP��N.�����A�8c�H�E�7W�������)V�M��1������T3��Y�du��3���+����������Y�9/b������ ������~7fv�t[��G����&U֧6���&�|ݘ?�|y
�ţI*f�M�A��]�*�S/J�7Q�	4��;rd�$h�;���$�ݐ�ۈ�|�ny֒C�.�Q��΁`�d]b/��6rB*V��?�3��zټ��U��g?���5�i$����^\(�EH�*�1�S�ʒ!�j6�5� ���,���A'�,��J��\=®���R��go�0��w'�\ͪ�*y/��,��0:�p$�M�@����Yf�D��,����'�@cIn�xվ!��Z���\�����ߚq�U���EA��v�}W3�Pd�v�������o��H�m[����H��.)=Z��@!C�樂Փ
�~y�;E?g���T�m^t�y�� W�����GG2�$D8u���&4���II�'�]�bƁ�N�m�?o���Ff�zcڈ�kS^�:4����d�9�Į�#���܆�1�	vQ��汹�p^�~D9��b�~F��> ��1��1߸܀E�?q���f�5��Ю�8��~��B�'�XZ�V��7�/+�q+[���k�:z�Gȷ���(��b��aj6�Š8� ��ht�ϲ����k�� u���mੳ!��$?ړ��~�,`��O��{�v�S藁��(�ɭ�W�*G�r�D��,'&�&��w����s"�=)��rW*�~_�g؏�#�gل͘��YJ��"��ڎ0��X����(S5U�4�9�왏��w*];}�����Y�����
��+~t�<�zW����ml��
��5�ϙ�F��J6� �z\-�\�X�Y�«XR����̰1Vsrx�*]�ʒ$��2)�og&s�J o� (o;i�F�%L3� %��]��/E�N7�.�Z~r�n�qKK-JUm|�oj�?�'�\_��"�J��~�v��C��o}��H����y7@V
��wfW.��h���C���[�,�:����N�L��;.,����#Y����B�T�q�g�X��!�al9fS8K*�4�.70.g=�
��-95��p���/�~�2�g���_�K>�
�]-�j��&�S����)]��4øX|��*]�2���\��Uv?Ǉ�ܢ|ЋJ�2uz�`ce��5w]l-��3\�^J�9�*d^λ�LƾYC���2/Ѕ�ғ��>�A#�:�Fd����|�ai�	�����G��z<�I*�./,��N���0v��_ҕŷݢl��}`�
i�f�LP]0�@�1s�oahWD�>�nB�>y�D��k�~vl\#Ѩ�y�ܚl?��<e4�|۽��-^�_�g�&�cH(*���T��	J��Yx���$)�]�l1��bT��Iu���d�f�r��19!�"DL�9�;2I7�(DSB�^�m�����U�{^��w�P��܎־[���{-�<���5N����?���^1/��e����-�k�$�����g;��eDTyj,�6/�2�)�Q�3&u�r��(��5��!ن}��5��3m��e�T��������qI?Z�{G7ۀ�NxA+=	���ź��.��wd:W}e`XP����i�f�D�H��{�ݕl-1j[Xݓ	lZ��z�e��pM��1�|�P�B~���l����}��������5��F[+��&%�����>�4��k�����K���w��'}��!?���to8�����bY����j�u��v5a'  <q��ݺ�#i@���_GB���ˉ:"iw���?�����q��k��o��ɛ��ce�ff|ecc�8����?��S'H����Ѩ"��f��0�}>f�xЕu���%�%3�79��c��Sa���dw���=iS�Q{�7&�W���(oq5,���XO�����p��UT]5��yr�Z�1Xl�=����th{]�z��)�ma�C�w%�҉��"�V�[�]��
��m�X��N��������84���c��O�M�(���B�mv�yb��&@�fٙCf�t���L�`���2q�����3��ȊW&y>��ܶ�f�]35O��%)��TJ@"�Q)ծ�ԯ}M��!��_$8��Yr�>~�0X���Q}��`fPJ�$���vF����U��i�ĻO1�!��ô����?wZ�ДDi��E�O����}n�󧴺�[7�V�a荘J�]gg]mx��?'r�'�&چ)�����8�"�J@�M���d�{�ئ��7@L�n*�5���ޣx��Z'�:�:�M&�є�*8�4�T���U�N���S�jN�eJͱ"��Q8�R��-X��i�A������6�v$��xǕ����y��H��e��?Ϣ�8 8g�	����)-��0P�j�  ���Ǜ�d�
3oK�z�Ƒu���DAd5u১�B���t�҇���o�KH�ۃjw|d+#�I51+���*��@�ȭ���n|S��ZBIw�gPdߓ^�-x���������������{q[{GIȽ�Rb��i}�>����?�h�b���bPJ�N��q��ٽK%{�_�P�(Lr�����ٴ�dh�K��a�0M����6���d2��]�� ]�_�4t_�fV�����ffb¼�(=Ǖ�-|�)Q�}yxqT�������$`�f1zL�硯2�( �hN4`)��!j�M8{Q9�ﳻl]��d]� ��:o�ui�!O¾��m�ݝX��F��({�C6\��Vh�	��87p�Z���5_6]���|_��y@�s�T]|�ɷ�	��<���\��h�\֗�2��e��Γ�qa��b�搩(�4֨VY����S�S?Ze(o�3��6#:���J��k��]I+k*�%u��$����̦�osB<�/�W@	i��}�P�[��O��Y7 �}p���TM�{�\T-�uZ-j#a�^�/[���T���۪`.	SR�B���T\-ZG:�����
E^���N/[�t�M=7�����:}L��vQ�r8)pX�
��h� �6u�ua�N�i=?�	�;�}�N�F
��J�q�],ql�R���k�9���El��$��k=*6�t8��;Ւ��h6�5!�5*�n����8��'��.��2'��`ҍ�u	:��+�%y�6%&�L���iJ
=�T��eu�_�jg����v0�Ex�����������ʚ`@D%hS.����̭ʌQtg�˾�.+o�
�H�Ң'�ZG�Ҭ�&�Y�2�ҞZ'�n��
ؚ��r>�����o)��US��r�u"���_����0&��n���ۡs`�Qc��TO�I��|�m�w��;�' �T^�f|�w�A!��&�(� f�;��b� ��_T�+�m��4���O$�����ga73�>}eYi��2��<d����İ�*�7sz��Y͚Bih��O�R���}��%�(cN���S���e��V���I�7Iy�^�����Aq�ʮUݣ
��\���m��{tČ#��"�.�!�@s[��-������Ys��^�K���,�0t�:� �l|(���<yP��� �+�
��A�o֪���ċ�N��U(��ћU-+��SExS����9 ��E ��u"š�Y\�w-ϸ�^���S�iD\[,��u�_�P��}�K��y.�T���q0�H�S�Iڮ��S_��91�j�z���4��W����RYb���z�Z�B���`��T�ht�=���� +�Ѹ�Cu�Y�.���z��&$��^յ]O����Պ!Cv�,���w�L	4����������8�n�sQ�)Q��������	*�b.�5��Ï�It5V7x���C��b�3ȝ@a�g	��\L�
����X����*�@���i_V/6��Z��A�<�''n��p}�VR޶�_KM+�6�S�3k矤���7��ӳ��g��{y����r(���x[r�o�6r4-*mp�ҙ�h�B��w�}D�c���o��0≞���E�U�k؎r���ӭc������)C���XH �I3ݟ��=����I�S��32�v�0=���e�=Z�-[�/)����l�Gb�����6�6������8&�Q���Fz�]�!�K�*6�&>�r�/�W��5�ܯ�k^��!���Y�]���2���4�E��s�q��
�˜?B��! ��_b s����[�-�&׻�6�e�:����R�"m�}�2;�V?�^��C���Nxx��ې�]9�v�A�����;� i�T�A��e�ר����⃱M8�������_�����	�:�4D���
/��E���q�x�(X��H���c52��~P�8'���M���78�>�@�e�FJ���XD��S�v�i��ё��!,�J��H�:WQ1��T�r}k=OV�F�߇]褱g����(z�H#g�uhQu��bgA��D(�]��q��Y�z��Ե�Y̨��B~���^�=? ������h�B�~/Qg{[�J�Ij��p"H>K�L�	�T�
hQ�\a�/�%� A-A���QKg�y#M����v�����k�	6��)b�n�!X �N!VO[�|4�JV����Y�<47Þ��?�!�)K�xJrC5� i���,+�q����N�VQ�����2
���';c|$��"t�u}��?Q��I�L�A�ӝ�jc1�
��� 2U��)D��*�����Y��d���~Ql���K��>�_�����Ī yc�Y}���vjȟ���X�<��{;���f���{�?�BC�
xz�7�ފU�{g����v8�]�Z��y�7�
����ϱE=��S�+ž�qΙO#��L�φ+��3�I��}ݺ_^�����D��P��3ӔM?^���>1��A١G�|��f����s��5`L,y�gS^��-�ס<���G������`��V�G�'�n��;O����]?;��5,z��{�D�
(0���+��*˕5^/F�g�0�#���XF@�ʋ�\�D,C�EqV��!�1�������$iT�C��� 	��E�a�e����Z.C�%)��x��C���������I�lnD�hf�ګ.Tg�z�Z�����?��m�<�s��,�\� ^���3��H�aME-N�C0V�_9�����B5&)_#�`���5UF����zF�8x\��V�o�T����~$c�o䍳�9��YEu�(ia���=؋֔�ο����t��A��ǃ�
i'�r)lT���)������`�?������w�wO;G�9���FEaC[ D�mOX�F��`{�6�:�ā�b���t�1�`����d��I��B����(6:VdY���?J#�'M�u�����J�k��ڹ9���*.AR��t<;��<��R���w7�Y��+�cx͗��;��W�ssݣZe�6��|E��HL��Hz{�;zF'o�>ӣ��qZ�f��~��I�Y"38V�!	5�~�T0`mt���~L$M����d96�)n�*��`��ϯ��[�܃��-8ʨ�,��9����*~���-�_=#a$���>��b���)t���L��U��e]�·��}T��U�2&��{�(hbʭ�Kapړ�d�D�1��"G����K?��q�[� ���܁ �!�/���6%3oFT1����=6�/��n��ᣱT#E��T>���A�q�~��yΡ�(�y�|��(ڛ%x�0�P��g=;a|%�!��[44��(��`��I6����n�0������4� @M��󯩣�r��A_�N�*��TBwA9���ՐՃWv��"���l��uP���T$�L���X�afIɿ������bpM!ݡB�yZB,hrS_���R�D��}���$�V�ԭc<��O]�#�²��6����Z�
�&oL}�'��wo	:i��w܆��%�W�$.��O�7�}c2����+��_����[�8�2�N��l�*F+����VK_�t���)4g��EB[i��0,Y��67��Ա�9���s�7;�G	��=C�}�!d7�n��OR�@�>�f�Dр�%	/DD���P>H���-cni�����O�c��j����	������F������#IIP��CL�����"F�;�!H_��
 dB��6�φ�^+�Sa|�bI �s_XW܁Dgo�m5f������%$��J	ͦ�~K�����?���]㩗d�k�Z�2�=�'^�I	!�BrW��W��/���k������V��� T44�}_µ^��]�T'5�_���⨷Q[�|~�)����^]�s���N�t�视�g�އ�{�E����POK��FY����C�@�OJ����/\bXj$�`�����bυ��I�}�)��{��M(5�Q�?-㟮8�m��M�O�(K����]�LF�祫�O�QeN�f�:�W��y��и�(��TU2��5iF�T���ͻ�*D�Y0��"�|�GRV��r����}��bJ������Rي}����z�	�a����2C+*D��lHǗ֡&��ñC2���GE��Zرy����Ci9�f���u�ma��N(�wZ<s��̿�9Y
�G���u�|�V��ۦ/K�0��G���r#nv7����R�%@=��U�l���v���0�_�"��i�&&��5���pg�$7�JC�0�̢�a%��7�>�(����b���OТ������ꝴ���O��YF�RO��ch��<�lZ�f�Q�>+�`�a���f`�������ڗ��MJ��-��߮��\��Ŧ�~�i�G~H
�n��=��A���\@m[��
6�ѩb�.?S:���}I��ߓ�����A�8�s��	�\��A��-�W��� ������������f�x<Š���7���Uw��fV����3��sc�	"�����AC�6��b7�ip�=︅ۺ>4���1�J�M����o��O>���Α�ڏ0����:�t��T���'�%�fg��y��lx����ۮ8�h��]�	�W���XJ&WuQu$��*bW�.ۣ�EB��Z�#*<�x�	A����!�^�+�,�~�x�����[���Bj�uY�|i�F�S�V9�BjC��ϊg�`�m*�]Ni��u� ���n������kP{�c��	���T�^�����X����P|]�<� 7�z�N��R&�y�B�":�! �)u��[�,��I�y�̨�����meheN{'w�5�ޣ/�;[�}��QSH�ƱZ�ۄ��F]Du����-`��f��X��w��=�Ѵ����y�֐tftl��сx/��gnW!����I�p�`#��:�7{sv���&�s�<&��r|Z.�GgBk��;
}#%�vk��������H
�5���fF�(w�:��w��B1��5�%�n����P4	8��{
��>1� 9�;s��W�����٣�q?c�3��o��C���p�׷o�tT�Z.��C��	D����LaM����Zf�"�U�����!3���NY��I��� D��8���ߕ�O�ro���y���l����V$��}���yv�Uհ1`��F`߀l���i"v�"�M�8i���ï���那�5�ʶ�4.���n�����$�{a����e�XE���]�.J���m/(�����K
e(,	��15��P�ɑ{֦	�Q�ݝ�2��9Iq+j�$���'���D8���x4���#\%��MZ>�^4;�8n$�e/�ٖ�R���+��s�U��J�ٟ�k�C�0q�#�4��^��&Y8׺�h�����k��=��&d�*H[>�o�ϻ!�o9cڙ4�ϡhF�R��0?Kr�a�(%�f�d�x!�M\�����X���@�jA��=���|�$���!�|�?>@^����;-ͅ�mX��p��6��&�b!^�2�}�N�c�"�K���##�8��c�{��jkqd��ߥ��'�3�%C	�����K�.I��W����'����n���C��1��	�Z��1�X�z���Vu���P���z����a )��sX��k�!���]h�P��
�*���kИ@���u�D&3��do����!0u�â_F��K
.X�o����ص���(|Ͳny˝G#+���2Q�� U�,Aߝ~нj{:�f�v}����>o��Q�|�j@���
�W��{G�K
�S4��)�ѵ�p�,�!5�#8�����jz�;�h��L �0��� �X�ra��&��zr/L��2Y�ݻ�23�Ly�Б�7 �w+0�
�D�f ����:>�����ι(?ŊL��?���n:���+���^+0>)1���)oqq���^��3fMF��� @���Y@`ˆpI��Ve0���h���|��w�%C�Һ��-R �s��v��d���}~c��R��)>��)�p ����*�>�mڬ�u�|l�$��d�������e��y�Ĭ�QuW��fH$��H�	)���+~S?���+�L�5���sv�8)Ζ9r��';-�����1��KkF/z��
V�[GP�終������/SYe��HCM�4�j���?�3�р����?\�$�U�1]�َ������ј+J�u]��AQ,٨�o���%��GԏLIԲ�%��0�Ƕ^��x1%�%����Zg&:�Ad]��E�]g�\B�����@�E�	�͑m�z>�jx_�з��$�#}u����!��
u���̮A�zel�&�fK���u�P3�	1�w[�X�����_�ǋ�]�V{����U�Z�鶤s��%a���_do��M�+��)�ӓ�i���f��]+�5��ˬtA�1�l�U-!&Lg�gv�d��~�d�_K46��*�b�A��v��\j?�΁�w�W[1)�9Ōߍ��j)��E�o�� ����Wښi��Z�;ج�&[7�ߕ s�+�X��)1	#�D�"�i�#�w�`��Gy�"B*ԗ3/��(��.�}�:qJ2�7�L��CNrQ�&&lxuޓ�	+V?mmB���'H�D�1N��V�ǡY/-v�]хZ���ћ�|��/[c;ƚ-�'::8n}��A;L�t=�Zc�Z�L]~ϓ�A~�I���r{�s��4���)�e��Ӓ��𥎊�FA���e4�ΤG�m�\��x���٬�5ߠ�r����E��D�*pB�5��j�2�i������;�<<��>�2��͸-$��\��+Fl������_
?��f2�lu�!8���囉��zSP�q婇:eK�0h�t��匯����Ci������eV���Y[��h
��	]K\x�z�Wjm�<��-���Ԩ8�X�����zC�"�}�����y����|FU3$!�	�@Ҡiǽy_+��q,͖�ݶF���]�s����f��
�2�
@���DA��W`���O�>��mkV�܍_���=�9< L�gK*���N.���� E��'`����plt$ ��B���4�6w�U)��m�?dҹ�4��B	�J�\}b$&;~�z�O�7T7C�ዸ���v�#�P1�����=%swY��d�F'��H�hl�-f�ߎ�&x�Gc�*E�dg̍v�1��7��r������Q�\����^�"�t�5f�"�}�1��2p��O�2���Zг�~��W�Ο5��Qg�.d��V��gQ��Y�-sׇ���y6UDA�2�ب��Ss���x���(�z����O�ٽ���b#2J���`���nl��Ki��Ʒi�QM�Lm!�,���l������)�ZM�Dy}����J����|�X �d��,]>���G^�NV j�wl�;�f3^+fHQ���F�xe�5J�E|�$V�9K���^2D�+U}�|��������ݥ��ÑsԹJ�ۤ�J�}~�O4���=~H
�9�#��;�,�D��Z��e���J�`j}%NH��s��,��G��eˑ��@��ۅ*�$L��fDY)�^�(}ے\��Ye�趐c�Wm���M@@h�ˍt2�S�0��Y���5�w�d����x9���`0Y��(qw�c4g!��E_*��@��q+�E�S��U�]��&n wl��N�-V���P]C�C��� ��&`��ZiAX9e�Ct��~�(�VC������+���y���r�k#Ù�A�v���
%�#AQ�~$�QJ9.X.��V�7�%B�_��P��P�.n�6�wH��]�N��n���������%�yGI�"�;[�d�D���8E=���]�6���!�������l�H��:��y�x���x�]z�XL��MZ��A4%G�`���!��۳H-6����r+�V`��X��f�����ਪ ��A2�o΂SL��A<��X�Rl�"x�8)^~A�g&-�Y񴟻��I{�lQ�ݣJL��@�-߻��E ��Zn��.�hL�{����,Gmh��a7�Ӓ��i0�Ab2�̿�Q�FO�? ��\�#����mKi��Êz�.��#����N�[l ����x� ���>�Z|��f�f���0a�\�-���	�?�'�yr��C�^2�c�OLW8����V� R�{������
��S���X�&.���%Fh%U`����A�yx�!j��'b�?@DU���ܳT �m�i>��8��gp=m6�]�jrA�����n�,Y��U�M+Fj��X�ܧ�0�C.I��Pa��aC�2	Sd���ȃ���c5YZ��@󨷥آ/�>�˓ٗ*����̝?Z�]�����Y�'��,��Q���~���/���}�k_�T��L���y����Ӣp�T:����?�p@�|��9�d�D�#� ���n}!�x0/����G���+���u{+�%��.�h�I,I׭��B�^���tR�Fn�c�h���wZP��O6P��n��� iu�Z :O#�ȺDN�3Y��g����N�7��u�b@܉ӚĜ�H��SɓӠQ�Ѽm��%�Z�����>���H����p��j�:'���N7�	I,����;O��ѽG���FNU���!�X�d�)��,�oC�A����/�iL�6[�҈�w}���0�H
ҹ��N�zR��O��������,T��\e���g|��=����8^e&N�����TX>����LŨ�� �X��-�p���|���g]�\0E���eDT� �F�l3|7��l���1.�V���R�&�E�Y#p�C�9�q��i�-��Ė�*�D)�0��P���
����Jy v\�֌l��ն�X�A��z����.�|��x�mY��r�΂�nZN̻R�e�
hdh7��06�nw|g4�=�X�W8O���c0Y�rҹ��'���Ƹ��B��(G4��w�"t0���5��lW��\i�$�c���w� �V�+���6���R��QUȁ.�͟�9vʧ�ݹɉ�?I��xdA�����gW�@���:P%�Ă tً�p�0��0�U�P���^�D�s�@��R�&��y�݆�=�^ZBh��g��xz�~���/N�x�Y���!�;�%Vad�굀8+���gaD�Pnd��{��Y����o��z>��.�/�h3�q��_脣2�[�KѼ��XzC,;���4��;�~T�/?PH�+�*K!�N�Q�K� �N�C5O`B��]���ĝ|���$������(%4� j�+�	���-r�
̼�0&��1-�	��uH��eѽ

Ф�M�	 sǨ��HJl��-
��/�|guIO�A�l o��_�!��g���Cw�v�Ďk���!.g��ip1���a��(�P���O�i��O�5�ǖ����CO�ױx%�hU�O<������}34�����A��>A�*���*B�S���W���f0��tZ�Y��	�Dtb�f0�t�@��Ƅc׎P#k�tw,N�Z��6�$�M���:~�B�ب���sB{�AK�����>Od��Ao��SVb�U+����졳���e�u�rk�&T��X�o|��:�4 z�Y��^��
�K��/��R(���Y#�bu�Xu'�����N�5Y�̉�����kܕ����`�9�R �@睓j#�-%�"�Ңu$S?�nXNGR|���6s��)xZ�EF0!�e�ҠK��j���y�B�����t�TD�C>N���#����,��"8��ֿ��X��w@�«_�m�+T���(ڊdh˳�����I��� ;<N�[���p�0��|��Bo��|;i�A�8��Qa�D�C��h�Z�̭� ln4Z��������׬r�'�h��l�J�:K��4
pFZ|ב� �G��(��7��6r�Z� ��b9�
iPV��px�����VN]}��ڬSE���lE�	[��䔀"�8�ȼjÃ�����R�^VՇ���JUbٸP����Ѵ%r�E`���Rz�"�{�V}?7)X+���.��S]^���^�Y��&��x�{��
�؁�������]�&�`�	^9U6�P�,ч���r�"n9�D�ո8V�W�rꤺD o9��S 1�$�Fjg���������$�<z����{���P�����:���,��3K:�@��NX���u���� Jdd�6K��ˇjJ���!N���C�`B����I�=��'�/W�F���S��Sg0-)g!G [J�G�aZjQ���C�h_%awٷ���B���k��L;�{I�;M��ܝ����V�u;��a�BY�e�t}�{M�f�L����N�[�j)��i�u%q?W�� ;���@9ϙ�k�|R6�ة���ix� 
�`����4i�6����Ic����l���Q{~=df�q�_�["6z��/�D�iEy���$Z����Ɍk�j$� Mt�ʃ�<f4�q�J >)���u����h��//[䞽��~5�;�G���v��i�Ě�ݷAJ�gx��]�i2���6�<��,m��*L^���
���k�b�����+Ӕ�7���\���	�f�Ϳ�`66}E�-�}�#ƾ��7����pd��E���P��}�V��\��ƫ��v������V/ d�̗���~�]�-�2j�'�p�*`;EuwW���q`��Nɒ=��+�t�"Hx!�� �_o~�M��_&��TGG�}�_�?�n1�N���3l��'��ӆ��Р�{#�B!h��|+�N�7�W�b��І_����ŧ��3���Ɂ;�J~��)r���L�_�8��sn��ޕ�3�t�濝}��X�3桳&(�T�>=/٤��!�^R��!X�r������!���7�]H�w��ye���\鈣��hN��HQ��C��^5�d�n�aY8������MXv��YV�Z��,���x�?/{[��[�Ϊ��y�0�m��p9�n��զXr���}Y��&��W�_�.�B*�E���(�B���."�r�m\�צ7(ހ�G2�I��M��9$U>��Vu��D��1�^�m咱��v̆՝ ��</l��蔻�`�#h\�[�S`��e�0t�!��-u���%Fj$-�g(.1���jV����t?�C���.�B�y�����kN\C�z�ܲ�\�� O���ѿ@�Q.�B��z������4}/��y~{�Q�_�$Lw�g��j�E��=;a������%�#(��|��q�TSZ�2O=6��@�ע�(	G�7���T 	�Q���L�WܦB� >�A���(�*�(c�_(ĄPL�mR����t�$���بy�*�m8���m��yR:<�H(�x�p�]a|Ĥƙ��:NDq����G��kjR����?+�~�O��+� ��2i��L��h���.U44��ai_!
�A?�o�*�f��wG6%�cs��]M�[��J���՟�R��vEM!� į����P�|6ȠI�
�g=�\s+��G��<x܏ぴ�w�%����YҐ�T\L8ʟ���d}(
r{��� �S�m;^֠I@	�y
�-���]aZ}�1\TWy���� �K��#�#�M!��q�m�ܴN��g�-w����o�9}
 �=���1�^�-���`g��ψ<�7zH�� �߱�*� �co~Y5�4+�<|~��G� ��$l�����Y>���ܹ7{�X"� D���j�\tKǫ2'� ��M��Z�h�|���%LL�*l��J���h�t�\�^��~Z��IC����q�B���*>�8�ܨuE��b���u�{�@�K��&����k�}��3�y�M�q�̪�:̿��QK�	��=��G��g��H���-������6����-�D����]����z�Ɇ.���c2DbK�+�pN����sK��M%2���5��s�c2�OW���*��7���7�V�iM9��b:!����Fd� ljeLXS�odo��_����Ŋ����$������!Ѻ���	���n/���Rcc�Rʋ�"�3�3�̘;/y�8����D"V����@!m^�V���%�o��f�'�(�wψ�ġϰ�L�F�6����a��-�t"Aq����HFk�����#�԰�H)z�G���T)�.�����'}^����8�V9"�h:A�$��9�ԣ����������x��1�@V�}hĔ��^\�U�q�p�;��k��q(iE��^9����t\'��Jőm�(PU:{B��D��X��dx.�^T��xF5bI��@Dx+%�&�()� aa��p���B���`���,LrR+�Tk��x�aA��u\S���Oj��lʇ�{Kc��:��c�$V�s����{�B>>�#���8����^��� �LF(�G:�K�}fG��Յ���S�ڸ=o��7����������4œ�����b0���\${aG�0M��#y_���H@+�uѱ�_���D���Q�C����Q吞t�q~�^|�]!��H��[��۲�1Bm��R��J�d�p�fff��zG�{�,��0Փ��g�ٴ�e��x9а��z�1Ie|���`rީ��T8TQ���n��XS�R+!m�� â�������d��:D�	C��bV�M���	�Z|\Y�v	�\����N[3[�oY�_XV�<��}�m��:�DI�:Q�L���\��н�V��$*z�	�ؽq�=}�i��B�I9��@�޹�g���XĢ��~�]庹�hAʨa�⟽"n�Լ~��n}���{���+���AڡW���b-��T�9I{� �����R�'�@��N�^V$Kϵd�z1��G�
��3Ļ	�ZO)��ȹzyz��o� 6J�b�&|��J�w�|�8�@c��io?R�=:����LFj������p���n3����2������%߭2���5��L��Ѝ�bQ+�v�0җ�-�ܰ�x��c%��s`6t���1���W-�F�+\W˩3\nz�S��I``I+0���,��x����x��!%�8_7Au����I��������:a���3],.V��\��l�����*N�7��\c2�D'��B�X�$+ꢃ�-e~�{���UYěs��R~8������K���Xu�? �ڙ�f&3�+�P�00�ڽ��|�� ".�4b8�P�F�:�UgN�4�w��+�	�:C�������rv�T��9^�rZ�7h-��#��s�=�e�V#e���������oц�2|�,��Gѷ}�g�͆��	W╪��Ϋ�C���ϡmzRلA�{�������sz���Ct�&�� ������{����Gz�k��.{q��᭶j�DJ#Q1�ŀ����9r�$Zov�z���5��q�B���l�����IPBV��mm1:w0BѤ�5$�� d�FTp�Q�����/�&*��ˁ���^��i�_b�>E^�}�ǁ5G��m�_�$%�c���n�	ͥYRYH/+�(��,�F�3��mmF�3�;����v�ڦJO5؅N�D~�2Pv�o��f������F�4�O��|����JJ����
u�;�`J/+5$"��x��[����z�ը��x� ϑY�5g�2V�%�#X�w1L�wjyW����3O�$5ż�+��Ǖ�}����@�̟#�"�����w�<�vUD&%g��\����i��!C&��S��Xg�ݕl6��>����0$<#S��}20a��%�:Ѱ1��ޮ��!���M"��ոx�S�#�,u��G^O^��k��H���q�!L�hgG��F(���@�P8�Kj���$���M��+x;Ufk*���1�#��Oz�	��P�HcZ�Ʃ��0�g0n�/�V����D0��g�u��?Z��kj"�& څ4��������jV�� "��U������'�kF��Xgf��xx�{�I�Z�\��h�{�v��Y�*���c��z��K-�4v����}����z4__C�L��1^<R�)�cL��,)$��I��ITBƯ�+�}ք A�<��p����qV[:-`�"�>W�dP�\��A���2!�)��}�(�@���.�N)EI��N�[qV��#�'+�������蟯�{�E���ا���?�DX���ǎOt��ņ��ff���7�k���.k뜗/ck)ЅN>��&�wy�������!C�4��f�fj�n�͞�����w�QC�Qa�rk葶Rh�?p��� �(ڨ�ho؇���B�+��䊮Y�H���S(h!4&áFO'nw�0�R[�����������\-���J�
������D��9b��>ä
_���H�8],��N36����b�Y2���$����^`�m�	6���e���!q��d��kL�2���7�Ж	����H��!_w�Q�I���𾾤�T,�Q�GA�_xW�cQ��,�G��p���w��H2�����܁³B<�?ԁ��*n�{���Hd�v�7#�=�N5l
�yvxl(�,�	�4>��������=�h�ǘ�k�AF]a_�P+�d���>�T*���$h'D
!�e�@�o�Ӿ��X���~a�	[���<.P���/[�����٣��GvڹT.�5w5�+�(�D����0�wTg���rz6�b��g H2Bl���M��.$D|2�����[���hW��`Ɣ=h�BPS����e��$��ai��H}y���h]9��C49�W�ԗ0"[*�����K�eMl����6нx�E���'��M����u�
�/|g�����!�Y]KZ��8�i���G��!*
/�F�:h-"�p2!��7�ǭ̌�I��>[�s"�0���J_����M�b<�6���Z���!�u�w���E`�s˖�%wIc�S�ۯp@�n�Q��Fe�|�,)��B��k�'l��@�I���c��(�Γ��\N?��
Q�mn����*=��=v��бk̷a�$��?Ν�Rư������vYx�' �A��]>�/�X���a���f��@��ۯyB�vgQS��$�$�g�^���WI�3C10�Ѵ�ZR<��L���b|�Ϛ���{:8K�HI�8�
�K/$���Aw�I��杅@�ⷜ��T/+[[��+����r�'����:��)�Lϵ�\�Y��LSvx�{}�3N��y����T'\`۹��9(��Z?�m�2-�:,@��A�=۱�5�-�5j"�x�^�~�dq����C.�'��s�q��##��=\�M��=�B��)�;��k���s��K���
*O
X_n�U(�2�4YJ���~��\��"�һ*��Y��0x�(�z�˲z5��Z#��w޲��W���ܬ���F��x
o�&N��u&~���|WQ-TJ�W�8����2�^&
{�3zR�&o�#�$�����OP�Ju'e�)�f�Z��K~�� �1U���^��+��Gů���DG��aOI�\�Kp�$?P��+��p�V$|�q�m�x5�"��f�3}9��nm��3�._���֘hG䒙�^�Z(����1�ZԹ�Y:̙�3x��͙��v��ª!��4�?�`v	7۟Z��/�{m�ݤ���#`�i�<�~�����Ŗ�#�I[%�O2������5;31�v�pKc%�	xg!BMZN��b;�6�2c�Ӣ��K���K��!�v?r#��t���f�S�(�u�!f�%�udy�"�a@�cω���$�+\ux�PS�h����t��� E��q��(98�����r��0΄|�C�dV*s���,mɑ��U�z�Xb�,+��g�s�c���9�&^����]�%�"�j�$,$ A�]8\�
vYR��_Y|[=Z�G��S"��Ȣ^��C��rBKgN�� �C�	�	,���E����>��U��bU"���<{��V����2ǫl��z�s=��,��(_�|�"�?�5>��D���yXNG����P>W!0��pн���I��
G�����,����U���\
G�F�X�������\4Y��Z�t\�F �Wq�{����H�XA�>�a�$e���'A�i�|蝎����W%=��	Y�|�lC�k7�&�~�ꆾϡ������r/L�"?��R�ERM�g���� %�p��6�|�ln��jEX���V�[wI ڣ1�����rW�J��D�ӔvS�1���]�x|�������N���֪�w��0��f�!ĲV��dd>6�$��G6�X������v'�
��z�N�������`[�%L!�:׻b<��?�v�@�8*�%9��4�1�T1��P��>mӜ��ή<��{�(���m �<N2k|�M��Eʳ�e�N���R;�Ϋez���j���q�
<���3�)J<Q�����K�Y��`\>^:�4F�M�t���/x���=Dz(#Uc9���gG�FuE��11��&���=Е�բ�K�e)>�N��;��Ͳ��k�u��wb�[���`[�p�CL�I>0q��\D�QƮ��<b���.X*�'�#��_�n�3�e$6	5���%ʝL�Ο�З�F2�ŀ�\0b��0J�η|DzG����O��I
�i���!/B�˔{ܔ�8��Jk-P%g��-�.��{e񉂃�8�Z�畸�R�$����ܣ�[���?+�l�����Op��0�	I+t�!�)�0�����Z\�:r�
��3Qc=��O�kF���1���0EqWqB�CP��D,���|Q��!j�ey����'�K����)-�H9���B���Fxz3�)��ݚ7��@��;u�hՑݗbv�Oh�=�#�9�R%��6�r6M\�%ya�y��{0�@W\$-�T���v��G��[�����H]� ɧh�ȷg_I�e�b_���zSU�h��Cѯ�T�%��bխR\��TC/vJ-Wq�r��#S};8
��ȧ}�҅��j1��񒍴��/���KCK�v��T�.�^�`t��_IJN��6��|g҃-��7�8����]'K��X0���:z"Ϙ���ľV��P���h�|0�+��� �=�m����8�c-�#�U8Z����@]�dk �.�)7�F$Ӻ�
��w��&u�O��"@Ľ(��F�	��oA-Л{�;Y�����nT=^	�Ob��'C��鐚u��8M}y�[��ڐ���[�@L2A��HW�@�[����L�c�F'���'.��J��VQ��НY2Vn��h������D
����dZ�*���0�����d.���pu{z����YX^��>�)��}��n��6%��ԅ��.��rR��XE�T|7i�>]=���`�s�vό L�	L^Uk#:��)
�양�;>��r^{f��u`:�D������$z�����m*�L�k�	\��@(�U!1j��<��!5p�Ιh&@)L m"{��m��&~+l�#����(�M�֠ʖ�<�xz�b�K��91���r	��XW��5Ə�o�SQ~���LJk9�-�Z��B��W��:����Be4�K~��Is
�7�y.��2kN�Y�
hO,��/�EG�� �Ձ���%�̧߰p�B0[�g!O_��x���ALݩW��js�B�� �R���@f��s�E������d��6H�jw��:�鍆�#Sm�ah�=�>fL~?�~B�����;y�#�x�ٙ�r��.ѿ�W՝jeϦ]@4�R7a3	���e�|�����X�XgD)=֔�8����Jz�-zGl%b���6����a��u���	چ8��i��u~��Ӆ�t�YFVj�׺J#�Cɕ
C��{G�à�-�ظ�޲ �����z�����i��P9�K�2�P�>�T�Fe�zW�8	�R��𔔼s ��u��Q��0 0�_�eY	�����N#�g1݆d�^Wv)������q�*(>�����F��ŲFhP���nwUCUn���ع6�N�`�G���ˁs��y��?�[�>�֊������2�d J�ϝ�1��B�Eށ�7����� ��N���ؤ��ޮ�����R�3��±���2��nj���W�V�����m�kC�O&E��_A���m�Њ9�pǞ�)*{���@5��4�
2qZ�}�?s��h�?���2���5�R:�/�%wZ����Y���*C�"@W�^��Q���w��ñ0!z��VA~�Q�)	U��6�M7�W�����U�VM�:ek59�B�b@�c���sǣ�Cʹ��`���^�Uֻ�R�x��)��aK��!�o�U�Aۧ���9��!�c	Te?EV=�)�^���[}�G[R͠�e�*��I��$�����I�P�KZ|~�h�.�tw��5)߾�5z��ֶWN�Ui��Y�hl>�NG��u%���
�}ro�+Z���˷�B���i��y�sQ璇 �{ �yN�n�����?%���>�pj(������A�Jv_��B�-���Wѽs��]\1�ԟܭ���:�������,��`K"�1g�E���Ҭ����2�Z1���PK��m�!�0�+K9�t��\��Y�XN���'|d���`��ԄQ`���!��	Ln��K0|�,�C�8��⽳��(�s����Z��#�O��}f��g��h(���r�o=�k���WN@��Ƥ��QbI��}[?v�+�|T�	^�,�t�J�����o�֤$6G"#�@B��~��$����I�Փ��]����r31�@0�`������<s�z^�[���ru(O��l��t-����z��xZ�4��{s_���O@������N�
6N��@��a��lcÆJYV%Wp�m�Aef�����3�v����	_7G���r���OY�׃�&&���𷬷i��t:�O�D-�V�x,��� ?��SX�uXչ�����Jau���(�/& Jn�ч�a4��y�SHC��3�)�#֑1�*W4L���q(�V;(�D�dr=z��A���k�y����q�q��-�8�t����QkR�C�`�$+�_�Z��HS��e���-���*�`&������6?��2��ܶǉm��o����0��"'�v� H4�w���-�!��X�����&�N%Ba�D���oI��x�8�KIh�����u�l��)m��H���l΍!��2��i|�E�6�5��Ƶ�r� 0��b`z���	���7�] ��iWd�(�d��w�6�G�q����fK��5�A������,��w�DL�[��tx�X����w-�z���C#�����?~&�[w6rE��CzßM 8���5��y�P~d��AKq3K�Z��%�� �}���&�@�
څ�p�\�=�gz��g�e��E�D�F��|�;ef:�N�	��ڎI��u����.D��{�ا�n?������7_���{��9J��EÇ]�D�T|��"�䜠�bA!۴���w�mMϧ�<�� ^�6�]��1��s�n)�����X�|�\�K&���S^�|��������3��[�A����*�9HA�!��w%v�o�-
ۈ�b�+��A��$��xv��N��vE�!�~{?L>������o|w�aZ����.�N�J���)�2��aGC���6��p�f���f�:���*I9 vD9x!NU���ܚ,���{��U5��3�}U-v����<q�~�K�_��. �������p�m_+&�V�B��N�fڑ�Mw���4(1�`B/�IZ���j�+��҈zH���H&֢��Ђ���m��2tu�G��N�zd;�l��*���"��YD���s�2�
�Ӳ��}�T�(�GZ`��G�\98*Mb_uo���G,/�U2�ᑒR�����?��7$j�� S)�<KyՕ�����swďD��zs�'��	I��B|�_z%=a����Xf]o ��%�6�I���}hQ��t��YR����pI*����0�=��7'~6�7D����溲��78��n����L2��O�b���4��;�l��yd�R��o�Wۺ�����{����'���QMn�V0Kk��]��-g�h	v�*�=qn�	���$�TҠ���=���z6�������O�<������E��v�Sn�?L8��yD�T�ᛙ{��q3�MR=U�Dh������)[�V:�Z!Ps��	Tq��g�!"�v��8��|L��G+�p�JeW���O�:�mPjb�� �q�HA�~P����G���|�ۄ�� p@W9ӷ ,���������WNK�b"E�OC���'�bC%8��'���<���9Dt!]��p���6/s��bX����rF�A6�'U]?s�� !�X�� ̙k��sX6N�	2m�3��n)�5�e�Ҙ+k��a�Ajy1R<�%	q�?E�o>�-�0����d6#
v�,^q;�
���<�9r]'�GA3����E���椂�%���O��łfOҋU�.��櫆�J��=^OVΉ�����/(���cg	x�2�|G���m��bD���0V��(��D��+$�d(�%�91��sv�(�_B����5�2`[��N��\��P�8�~�_�A]���a|Y�K�+�V�!�����Q���B=����3[�$��Z�}Q��U�pe�u ��{T��[�a֟����R���-��_�z� �ݼPD�D�����"J���cY�����U/�/3��'�����'GϺ&��l�gw �3l��٥�D�v�}gT��[a�Y���"`�|t�*:�vA� �$�1>�d>�$��e	����)J�rD�Osωp}�=_8��������6$t�T`�
��4%~(�Y���i�`��q�0�b�'��0c��+l�L,'�ъM�������;'+[^4L�4�~X�n$��|�Z��C�J ;�l�sX�r�W���L���c޵WՅ�rM|�
-Z�\$Go\�.��BD�O��s��i��fQ��6����ׯ���7�����O�흻�L
�ɒmȺZ=�s�q�!W�
s�?u������_�N�r,� ���r��ke���2�G� h�N�
�Q+��c���kEY�����V?�q��$�����!���uo!��B=�����Ӝy���HJfn��x�L]�j���.&\��9�ڒ��q�DFsj�S
�=�`Xr�-P�vJ��b!���҉mj�b'@�3ȵ���X<,ǆ:I�3Q�p���/�C��W{9����+�?�}�l���	�B]��a�>e��P���jɞ�é$0���y呱��&��ﹼ��]p���7�<b�p����B��yS��K�\h��+Y�#�$��T*�>��yH`�7��E����e��gD5��z*1��O =f�k�E�����8�O�Md86e��	���q���/���,S(∾h��p�M_��{��昳�rʭn� L��ۨ%���¿�ZD��!�k/}�5��4,�J�y�otw���\V�o�N6,5�'	�~����Y��E�Γ���o��
ch���w�A ,У�˳�k���Z�w܏#˹�K���w�ᔶLi��@Ҕ\H�����~&��-[�z���C�S�փ���U��J�W.�G�l�)�*�V�1Ւ�E�r��y/g'��-�wQ�"Ls�ބ�����^|r���ԣ���d�� �D���$�琔��U�W��̎�$����ڼ�T^�e��FEP44�p(�T�������(t�]7Z��2U�\��M~��C+N\>��Q�3��g�\?�NŶ���;#�~⠒#n=H%�tB��a��f�+�U��>Y	y���Y*�\[X	˳R����=�7g�E�Ѐ����-�+�����|9��E�_���n��8`r��~wː�a��%
#�"��q}��'*��TG����(]3c�)�Z�F1gH�����$(�{�:��p�4(����5����{+/]�r�*F�5��C�}��Vd���,��7+LL�������;���,4$΅?'z�<������7ݠ�Y�1�\JM��W��~R��4B��y�=	��8=)&��V�>Rm� �&n@�Gd����_EA�s?�`��`�Af)�x�=�����$�-n��򏪜w���3^t����[���&�F�2�L�9UN`Zt�[��c��o�חU���EfV�\��� &��i��I�^|I��p�Nk������MY�˞{���3��}\O��J9c�Zߛ�������1u������:|���ĔJx�1�� 2�w�E�^�q�vU�ti��,��s{���mg����Ǐ���=��fv���nj�0��m�=r����e9$
�3i�=�J���.��NC�b(-��~j�G�5��X�ޯ��,������H�ju�j�R�P%P�,< ��3�4��{�|nZ�s��~T�H���Jbw�j	{<$->�$nG���Vqja��B�2Gk/�X �㸠��~H�	��V�<; �n&�� H!���jU�4X˯�jm,41��`� �{ߙ�= �hՊ\q��%�!������	 p4X���g�ECF�c0�[���;�� �6�}����dK q��UpxQ;�03��-�D.�uהLK�O�y�y�i��DO�
뭖��s�� ����E:��;��u)@U���c�o���?��dYy;l�!��S��Xl�>H�'�%�]��5�]���S)@�%�g�_4��	ٽ��%�M"�y���w��� b���{�z׹j��8{\����|4Of�qaK�|������R��lary0q�y��,�j��?�e�ɗ��i�`}�!��+z���		�?�l�EY��M�4���؃ZNq�W��x-!RW6id&�u���Ge�SOq0CtZ��E��;��$^�)��O;�yT�m�:E���v�ь������f��}pA�j��.
u3Cfaܒu4*�YJ�^�����]�a��f�M-�'�sfET�i�P9��l|L?����5ذ�(ٷ�ˈe�~:q)	Z�o�u�̟8��^��j�	�酃7�MpN���k���Ɉ��>�|�U?�7�9��%�����rPR� H����j( ���D{���,�l�B�,N�{aI�2�%�q$\�W���H�S�3��P�N���N	��	[�]�2ZM��uQ�4x �Y�9�ԏ3UY#��,�Ӵ��</��Z�8��Kk)�qe�1~��+�{:���!�17���t�H����l�L�-���w��(���FG�F��V�P�&�\��֫ ImL"GEy�����s�+h,�m޶��lV���]���qcV���0e�T@x�'0a��-�$A�ǙE� ��Gb�Z[�<�5�L� +)^���>�b�Vn�LL=���~q�{b�K�cO�Z��C�@<(m��u�Et����m0����?���0�d�,/�d�I}3� Шm+�]�~l2���08I��}�T�`Zǌ)l�^��M����fM�&��$�I`t���ƻ8��$�E�(��۟;OᕵJ�ɧ��2��	����v�P|wg��Y��>�|�~=�ᣟ��i�Kפ��9��y�w�����RcS����#�[L�d���Zt�]$�>�㊳V]�$U�:Le�(_����x�X��S�0Po:/�A�YULķ�L�ҡ�Oj�)���)N����)J�k�^�f�Ü�(���L�;����[������`P����!��LعN��lmJ���/Op�M�<��Č�\]�~��3���֨5c��axl�
�u��p���Ň��h�s��F��"�όjX�;�cj%�F5�����|d����p���Kid��Vgјc�����lNp>pn���M��+�t����������,k���2G���v�)%��� W�%�W�z1ˡ�+~��l�_3:����/ wณ�{)����/a�H���W��8��;� ��S����LI��LW��0��SK4��%$`��P�`��s U�`Z�;��z����-��VE�K-����2;I����ԍ���זJ�1��K������6Lۻ�9+�������4��Z]T�qz�����)�7ڿ��	IKZ��^"��E��"��?�z%�-6��%�@��=
�¡�H��=�Ġ��乤�~�%�7��N�Ϙ�)-��<��5Ah�%�*Xxȁ\s�ͣ/*\v������\�~��lʾ�Mq�����'
��	_��T)�C��u?��n���"C�J��m"�Ki ��H��g����/��Yp���e5TN�-4���S����f��t�V �TH�a#.��x�\�^B��䦿H�ʄg&��gO�C��p��g�N��4W�6��^�ȵ�Y��lC�H�_�WJ0# jD7T��_��q@�#�i,�.�W.�ȄhX������g�{���ڒ�S��1��� |y�؋�xؘϿP,�*�VۦKe���Z6�v��8'E�@�ܓDzx9��=�;g
n;��"��*ҴRtQ/�����'"b��^��Z�߭�
���d�c���57O�}_җơ���#H�K01���;�ۀf�7V��T�^ӜJ���VT���wzR<M�63��ߊ�]x��5��S��Nsˮ;�LJV���H�A��F��]���$R��K:�=/�f��ts\*��v�'�L9�d��z��gU�Ģt3]��,>�kԥ�p/O�,�d��*�s���v�ڲw��ג�����L;O
A�l��1�.!�{(���R<�������I��8�lܹ٤e<��ڹ`5��g�*�����S�C�R--��II����� |��l�c���-�1Y��b����ŵt��p\�}�c,�L�2�������rƖ��p��|��]ڞ��� B��9�$��m�f�n&��t������������*�@q��3Ƀ)�g-���:=r���N���M\'.��[nk��f�7A#���<��Q�[����b�z9;�j��f,�e���|d)Pzc�?�+.H0
5�_�v�O���\ֵ^��v[��lx�@�M4J7eC�`��a�z)��\O�_\{���Qe��a3�zk}'����g��~�DZ�N�fd}j_��g�BHU>�#z�Y-Q���G��sTx�	t�D�^�]��i� Eǃ�[`_�H�X+_L�o���k(���ہ���n�ʧ�I��L���u�Ȉ�F���#��69tX�R�1��w�L�v������!Y���,�H\�9�{H㬸>mc�<:ǩ��&�_+��L�P
��q�.N{w��n���E�o��.�+�Ed��q���s�V���p\�'�:1I��������o'�ԛ�펪Z�Sc`��4����f�h�[c�bB�{���
���p������S��\R��9��7C
:@�׽V�VC��,(F���-aϭ{�]y*\S~]�xN���!p���& ^�_���?�v�LW�hQ��7���alSb?i�����w���>�`&�_���/�8��p��iD1^�8�\�(�?�/ޛ�!"��_��k��P��c͓���B�-����l�A�yW�&H�)��4�߸{��Y�/�a�e��������}r���&��ަeܞ��L�g4��B�H���e2����	R�#{���(p�s'k
*�D9sp�Vb��q�:�bF �~=�c�05�� ��q�E�	k�ؕ�kЕ5�#�4;!�>c��x�� ���Ü-!�h�E8�G�������]7n��gLLz�w1 f�0?�I����Z�K���;���C$}L�{L���O�Hu3�	��+2��QM�_Z϶���g��ﹴ��U	�cB�ֵ�@�MVv���.�u���|�0c�R�FwA��4[���Ak�F�'�b�O2�_�㉳��3}��������,Ӹ�����!(&�U��?�䆐��)N�7_��.������s�Jؕ���B�Va6���@�Pּ��r���O�I�;�1�Y���Dy���Y�E���<E~&�;4(˦P�'{)[�K��֨�j���e��S����l��ߑ�x��20֑�A�#&�$��l4!���#���Zp8�Iq����p7�]}�����~b��(��
�ݒ[$���	54>F���qCk��^�����ݯ�,�Y9�u����C��z��R��X�nz&2�D�c}~�]�i��B��V��t�O&��cNV逛�0Cr���܋���K׉^�l𨁟���w����z�+��W�5���:l%�x�
b3���q�B��B�5U^�Q����L����$0,,n�+;���d!���AtS������I������;��ԯ��}/O�-��M��%��VVө*�:�H�-0�,R�S���n�H��e���1�E,!�n�[�V*(��Y�n��Уq����T���ICɵ����; ���o�� �Iz�?^��Z��x8�{E�F�z�nρ��̙�5����`����kA���y�@ԩ���lC��.��+��+f\���pY?;b
�#�q��#�����Q��\���=��+�]��!S�)FC0@Tl���,/r=ܜ�1J��e8h�r�������8N���<��ݕ.��OJH����.T��3����&�{�z�����^$A�����rm*+$��3��3�e��)�Q6��e�#A~3�qRV�t�C�آ>JM�w�:糏�j�|Z�]�p����"���'-��;��_w�=�x�.N(&^X̔��q�`���cg�ߨJS#���*ΔLjJn�`R��~�S�3X�,ߣ��PIP�K~~����d����<� [�u��XT���_(�����"l���1h���Ux��9%TJ3��vf� ���-I��ω}Z��b��T8t�g;�c繇����ܿ�|!�}����Kϻ>�&�����8�˛�1�`��O�Ǝ��ڤ�U�
�J���W�N`I꒖(�y�����%ʓp��D�D���BD�<�����m�����"=�����Ș�[��Y
�$z����0:l���v��Lxؘ:�`c��1hv%���ފm9 Y]�p��p���:��Ƥ���oD`;˖��)A��c�mUfn"�Z��>��˽?���0�q��Vj��{/�Q�������~�#�A`�Q����"gjNQ���4�:U^J�M��v���>1=�Gf�lJI*�N�|v�C���'�hf�O=븉���r�aZ�"km�dD
��8��v�L�.�p�i�-�.? �P�E��#ܻ��cG)�\[_�"z>�(��:��P���_Z^X4W�hT�ڒ֦��=[��=@o=t���������-��l�Y���L�q>��v{i֝��S�s�f���������~��7���/�:`�w��R~7���A��h��A�)�Z��I��t��b�;:,.��lFL��a���`��$w�"s٢#f��.���3PB�.����rm��PGb����l���L�/���h���h]���=���.*U���j�z�h|"�E~s���c��F#��c������89|�Q�J
a�b�(�rV?���a��r���0��*�͏��J��T+~܊Ʃ���FS����Q�r��6	�iG�����6e�Ѯ%!.yw!��>����U��PRШv�t�i���t֭/��HI�o��7��]:6��t����L�������27�z�w8<���wW(�� J�8� �6�BW"����|�:%�d�:	g��G����y�R�?���|�爆��o�&�Ccz�-UJɬ���i'� �$�6>�}SYa�`��Lq�'o��|�#Wζ^1_]��ƺ!��?���EN��`������P,�����R��q��ł�u}��h�u�N��<�	����h}ǙѼj�f0�H�IL[�M4z��<��U��b���������ʞ����s`I��c��e���g=�%X�n�D��~�\ŽUo�k�f��Z	6��hv"`�JMx�Lb���c�ym� n��PrR�,s�:_�'[Rkx�/��.�p��Iݧ.x3;�W��9���������ɱ<�h	S9��-�����l�m�M����2��sn��iF�
=�����F��*�n��e�1M|�TZ"�#�6w[؆ ,��P�U��Dڀ�'�ı{�D%#��r�|a��HD����}£&ˤ�p�O�y�l{��ad�K��DZ�|'�^=Ǩ�h}�P�`����ҧ������밝���w&PJ�\�!�q�|�7����S��V���⇧fwfQC�	�=�C�۶��~��4]�e'b'>���j�m7%�o\�ms8����ޔ4��J�*�5��P�m�ī'���9�N)Y(���`#�玎�o>ն]��a�'3�VXގm��"�\
�2���B�/VSq���,�uy����L`��WIS�b�%Ά�E�1�EU��̬��g5�"��cN��X2��v}lD�g�"n�!��W��W��睨��#1?U`�`ps��<}�٢��fz莶 	(n��Ӥ�f�g��aZ��m�j�{<!���<G���X��A�f���R	��*ľ&�9=d�{�қ����ր^������l>�C�_L&(��%�!t�1u}[�s�W��xW��n~�(|����zW���!.�a���B��r��S��w�g��3�XI�4���<w�M�U	����\_�6��	1�:���C�F�oF��[� �8�ڵ���sn�l��]��N�iʋ��
�L,Db?{.�����,j�+w�\k�����dK������9-ɩ���`��I����xtl$��3ٯ�R����)w����΄�T��Ĵ߅�`!z�?꒵��وvA��x��'/ u�C�#��g
�l�o�_��� b)�q `�&�+�k�I ��&j'l�d�Tܟ$+A< L�^�Top}�j�\�Ғ��N�5���o�������&�CN)+����BV���qZ�!�d�w.i�3Y��l3���l[5L@�Y�'d���-�J+�2��]�!v�/��� �Y�4!��.Y"��f8��r� o�ʰbFY�y=U��_��*����Wc~R��7���CR����A.�|7��K�|f�6�K�B��!J��Na1dt9�觳!���t����X�骣>���}�+�L�r/�ȡv�/�r_�=�n�
��Sߢͤ}?#�y��N����yn�z�7}����yk�t�����e�#?��8o�p������.�����\|T�}���:�(�F_�v_-[v�v|�0�k}��F�>��!��=C������j����칔ߺ�TME�x|l�s�w|�K�u�UϚxw#�m<�y�Nj��fj�-AhXv��5\�����]/%r�W���
���%��N�rNkͥߨ3�	2���Ĕ����PNI_c$YDd�0�TM�+����m�m�˺\�GT��`�>�R��e̋���V%U���+�(��վ��a�QɄ��Z	��J�K�>*�qD���j�h����C4S�Ws2�YK*A;K����?݃�i͢Z���K0�t�����􉃝�HI0��y��Pe!�����!o�,���>Ph�w�i6瞙*��(��/|M]�1�YM<�P���׹�Y�����6���X4��a���Q�D���������@f�l��kK ���;H�-4�f*s<����B�<�p�Y;�Q� ]�_��J����x�2&�������0��7��Tܥ���J��
�0:[}Vo�dƆc�O��b�5���N�,�D�u��5Έ���|f0>�o�P�W-���:�@�e��#Cϟ�OD�����C�?Q�k*��~�r�q����4�h�L�KJ����{JM�F�1�|��xu�=�^���[-�c���ح��=�V�O���M�+�ꗕod���~WP~`��>C"S<Ԡt�5��]��5��Gd͔��7c�	�,Y}A� ̖A*�j�Y�s �ki�mLNW�M�~Fv��*�pqלхt�Tu��yY٧(�"q���A?�ۘ��h�S/��|�luˆ(!�d���IG��r�`����e��ܝ���8S~�����Nj_!�6�������}�������Eߛ)����DD!�z���:_c]/�_l�$c�[�,]�m�kY�{����$���j�3`E�`U�C1�c��;A76�l��
�������#-ڬ�xb�
ڞXW��f�(fg�)��Hυ���Ȗ���;�����y쯵Q�����;)������V���zG�sidZ/[&�n|�H��|�ꪓ}D��J4�1��R��� !�Ɉ�&���@�,�49 ����[�"�,���v^�mr��r�:��|�K��!Hz>�
��QN4�&��Љ���0�V�P�b�?�dՁI�Ȩ?�ڦ���Y���:�n��F�!���I�C8��Y�n�2z4�Tq	�h��t@
���� ���yep�����Ζl��!/{��L�y�8��8�|&FD�|�JwfQv��_^���"{Ź,C�W|"���=Naۘ
= FCv4�đ�4.��!��Sޔ�9�� ��o�čk���3o�D��!_g�����iv�0�Y�'P��%�ng�E))��s��/d��f�����=��9�U�i#A>�j^�#27л?���C&�y��0���$8 ���)�v�������3�*���3>lwH�ռJO�k&��<<G)%#/ưcb����'_(�3ֹ�S�ظ�$�`<�x��\��~��d:)��Ndl� D�0�R�f��;n7
�Ϫ������x����3[mv2(/:���A NjJ���>���AJ�,�݇
o�ي��]�t3��v4*΃���_ �8ϬM?ɠ	�:�(ޓ�k��G�,^26.iK���\������v?����Kܖ�B�۽�]�F�� _}{
������r�a^����F��W}a�n�9Q+��زXP�a���H�ԩ��_�V$6��X�T�c0o)^�I�ʾ�nu����6�M4~:_͖�"-�>lC�������Mz�%HtY�B *q�|��N�V>е�b����lZh�s�����u��|�ƾ���*�#���[|P��@�9V�;aG�W���!�&`�pf���1eK)�a��4U�r�#C�3[�]��p��_��OH�Z�eŤ\q3�t���z��t���X�R5��=�PW�v�O��`�e:n�(O�gc�֬Ax3rޤAg��4wG�����z5�d�S�?Z���.�"�s)|J�$�{�\���i}ӡ�LC��d����,��Ny_�Dw��-}�z2�r�;?�%ÞuQ?�cG�ֻ�Үzp����*��P�{��g:���8���!�q�g��ƶo&{AӋ0��ܪ��Եj[���>�A��9F�P�G@��!UF��S��S���,ۻ3?�ǏF:)��X���V����x W ��6���2d�{�=m���cq���"l�;l�2�T�e5i�I>px<��tL�"��_\Z��ez�R�������%!\�Ci���}�B��l��tG��q��VR��\z�lGu��;�hњL��k���}F{H�H)�~̀ӊ�,�⁴���z�Rk��{` ۼ��v��[�,�5ń�H>6������+=H�Tb�ӢO�9����s(����Rx5�%K�K@/mB��q��W7�	�/��I]�$���Q?�$l2�G�(.p_��f9�5*�{���I�CQ e��F�|Tk�6�!�D��*�x����1��S��2V4�|��B��&[p��)�Я�K\��M���T>�%�~ʡɀ ^)�9P�S�d.J��v�������7°�)+��`�ѓ����0ܣ���~ $iX���EW^������G��2 w�X��zσo�͎�$�8`��n���HZ8C��������)���T�\ߏ�$:(�2,v���`z�:��obg ���C?T����r�vo�ѓ�X^(=b���qUYa�JA�/�*��#*�W%:/����9�gЯ�F.�%q����?��<f�����x����tS<�.6o��U�[�7]6�T%�;Lc_�����I���n�z��ϲ�x��6yj����;$��Hn�2g$���0O��*ٌ�1��2����ޏ@�KʏO�U!��p.lWvS��|^L�bh�3�f����7y�4��i���m�]�p�Î�K�{�}%.'�~����&��5a$�O��>�2%۬����A�̊,I����P��]̹���^{�#�f=+|�]�P�"h���<8݇�R5��*�C�B�����pd����Yg�O��+�T4�SD�]�5�����/&!-ս������\�X�#�����=|6:�S/SPG�\tY������sK^�O�Z�`�PTC�ʑ���9��/��Ǝ"����*e��.y]�1&��o����;M�$�Z�U�A����z��C�|V֟D��.� ��a�TW�1j�z*�EYc:���H��)o�~m� v錯I�%$}E�QD!˘�žji9��O>�\Y$k�	BȠ���ǔB͘��L�[1w8��P���*PH1�!-C���ۑ1
on�zuO��N��^#��YT�ɖ�"/Ce���Q#����>Ob�&�?Ƹ����A�H�ԗ�'/&l0���M�ե�|����L���D�&����^�^ m�Փ�{��z�����b&Z��+V?����	o\�,�&[5����OZ�n�L�~�G:A��}q�Ǧ�b�厔�St5&H�p�'
�O<��f�j����W[�%�7+g��U3N^Tf�p��I���y����Rg |��H��w��૳P���EJ����t����e��&BԆ����+X�۷�hg��G#��5s�b�z�����G����w���;�e��+)��V��I�1����џ�6Rjbl��8;��9�[�.�a/����X{����?$"Qx��HßPXN���c-��>0�R1cn[(��& �t����@Z?�}���is&w�3���_Qx���'QKK���&EZ���>}��J�8=�B��(uXx�o�z~ʢ���Z�p;�3����� D2���z�������BM(|�q�����,�L}���H,l�tC�+G��,0�p���=�z18��i��~�� �Vڂ�����we4:�JżOB�[N�\@�~y�P��J=��QD2nݙ���� ��K{����5�	��������_,tn�g�Bs0D�I����D.���:�"J�<+��f�T�`e�@�sV1�Q6f�*��V�BFN���gP�!�v�9�,	8����N!z��.�z�3�kHQ���$� )����G=�m(4儗�W� ��_vV�Dz��N^0˸y��i�xM���!��<~�^��1�� <�8�M�;���;XS!�p�;��{01���&@�4��y,��R�������<m������3
Gԣ��{R�rNC2���S6R����ns��#�+2���\[ ���.����e����9�q��פk���ٕiY߻8�O}���^�'�yk�����7ɇ_�c#����)a~@�#���c���(��s�3���/����H��jB�n���&���$��]��8ć�Gw���v�	��%C�{~y%,�1� �l� �����|"ݚ�^�]����Jϝ�)֓o�'�d5F#mMp6��M[~�i�niH�By��-j7�I���$z��%��-�"���9!�h�<�w`C��I�8ͭ?�[�jTL�H�g�E<�D�������Ƣ�}�!T9��29D�N1wZ���&��ͳ��n8I̬f+ƕ|;@ *).)�7��u4 s~��̻�6����L�:~G�i6�8�˒[  ����A}]�aIZ�?��6�NJd���M筪tE��6������mf�nݗ,
���Z��@��!����,��	��/��Cr�C�=�%v��ר�M�����ܷ�2� /Nߤ��ǳ��qn��Z|��'���+=BO�eϴ�`s��fV.<� �~����Ī)d����S�)�8>�
5�D�7��MS��xE�u��G'[��:yg4,k���y��P�:���܉
|�����V���np�͖�X��dس�U�Fwhi�u���P�X�A�ϖ�?a��	����5s���7��)Ü
�a�X��Q�^N�n-�tJRɊ� ��v�7<^��&�D.�9�S-\�t�a�]�ԟ�]w�u*��r��ϲ� �@��}J�@�k1zU�SΧ&!�i �G�B;��փ�����;�����xvƞ�X���r�-��T�����i�l�����4�
%����AJG&����jq�r/���/,!P>��e6j�,�YD���K�r�	SaǲTK��%�c_������L�2�v�Z05�s?����I����y:#?I|���iY� /��"M�6Ms�ƣ�n�;�94�n틳,�^�D~C���$A���W���
�'ɕ���R�֊�RNl�n]��w��6R� b0_�-�L?�c�!��W-��yv9pT/)���^2ct��H����Q'9=y�fIw�C�e��; �!��xv��iբ��\��75Ꙟ����3� 9#����ON&�2d}�&�6M'��(�ғ��1{������)�N�7�.,6?�*�& /#�:M��Þ���ͺ6�\����N��S 2���$�߬�竛�����v���w ��\��qH��:��4�����ۭ �f�mh��&�. P��w�X�P�r8O����sF�ɾ��0\S|����v{:λ��X;�qcl����f��Ԭp���Q��Ό�X8{���/�f'eu���Ɂ�$�Ͳf��9eb,nS@['u,>z����L�vC�X��4@�2Q0s9�%"q,x!{�H? �%�����!����k|\w��u[P�;�S@_G.juP8l��E�}���x�G/���2Ժ~Qtf���I����Kھ/���{\Y%��]%���3�v��p`"�K��W|�9J#Mrd$�SD2I���kO61<��p&I~�f�@Y�K�䌱�|�|����"�s�M���?#2�����:؎qq�#�ꃮ�3�$���[3q�������������dBhw9o~Q�) z���_5��Y��p9E:|is3l^��~��{��<dN5E�	.�H�=���蒐�qH���K['�Iv�k��,�3�L[c��[4u��n\�5�gA���n5���bM���+��-�r瞫a�Rz�P.�1�c*�م(w�QiR�14��z5��l^G���Ѿ�x�T����c�_���\6��60F�b�`�C,��c����v���G�g.���r����>$��R]��l�;���1"�Dt0&����$]�����8��|����K�W�P3y�a�G<_�������Hu�+&dѐºeCn~&��3�ٗ�O�N-�YL���%8a$+h��*ń�C��ɉ6�&g�:��[+��7�/>)���dm�=��wO��7U����z{̆7@EU)���
㬉Q;�I�Y����'�[�0�J����ϭbׂ��D�%��n�(���u��c�q7I�����<�Бv�&���jsՋlK��7��'H]�W7�2��"_�L����S�����8J�`Bs��q"��������&w��$�y-�$4���;M��"3�Y��s������m�FW�r9@�i 0����yI���J�x�:g�L�5��0�}�p���B��/����$l/ݟޡ�OۃqA�D��Â<�7��M����_F�n���_��ZO꬜�uHT���0��q�HL&!�A��N�J=�㶮2�{���W4p]˗u���2����5�3�g�!po�ZwfxH�q��n?	����ԋ�.�Y'�����u�i^�-|�T���;2��\�;_�����:���I`ot���@<�B�3v�hÄ���)�Dd4��0������N�a�i�P��t��'��G:����ރ^X�A6=��ԧs��{m���gcP���]:�����%�>8�qS�$���cU���e'5��հ�9��,�4�׼�W[+��^˾q|��7���ў�����.	�v�%��ֲO5������$a������~��4މ�?>��]k{@�����a\�ƞ8FGZ#o�Ԅ0.XV��)��3ZF�Vm��w���+�&��+����"��g�K�b:Ҕq@��f�mqGV��}�� ��̙���oD6$�7�г�S�wb�E�s�H�Yѹ�05�v�:����� �'Ҟ#��t�{[��N��_aM�����)V�C�G�9�=�&�Q��e`�����%)�ta$��B�G�Q�.�0�Sm������0�C2�5wG��({ia\g U�"��4�u1�V�JU�'�Y�خbn�Թ�������*���A����W���.�8��d�����k�)Cx�n�=F�ɦ+�F:Q�4��� �j���un�#-S .I����@�l�GS��B���4� �$��`�;�)��}�pԊ�#��y���bq��i���!rɬ��n���T��_I�.ގkA��h�0���+x�0i���y�R�$C��ϋ����.��i�qE��F���7��ɐ���D��Y�L�vi���/�~Dg޽��M����{�V�V2�d�E�K�.8dX'�n�e�>5�R�"�3�"��6s�+Ini��s"���f�Aʓﮠ���_%����k�"����1�Y�I�����kU0�&*�К��h`�(��aH&����x<[��і��t��I�!���x�ɾ�f�LK�$;;�AK�0��L��U����&�7�L:L8��̨���q������,z��V+�镱��U�B	ZbWfh[T�&��<FH7��9��*n�X-�9��8F�/�c9f)O��I��Aj�e�=��?Bv���@�,�l�Qt��յ)9�P�v���Em;�e��'�:�W\�Am���p-c�s^�����=� ��������F(�=�%'-�7:S��W�)T
.�/�>���L�ErsL^�@(%�bԇ��bL���E�xފ7�4�X��3���Y;�]��{sOHa�nyC��m)TY=[:�`�\\�>]ʒ�L�^:}��A�j @u)��B̙<M����F?g^V�v�6xx�&��� �B.if)]�w�����jɶ� �J�*�bz����]�m��/g��]���\	����?8��+nS%C�qqJ�8��fw�����RTt(]�?'A�J�ȵ-��EP=��l��_QO�߀�3
�{�Ko���v�m���tX�BH?�At��1��\�������$/g#3�x�#�]m(j�](��e'�W�*�]R�?	����G�Eaɯ_�t�s#q��(���m�k�h~a	-�A�������f�H p�`OOoX+V�*dl�Xf�7GsO��&(��DM��]�\�j:�T�a�55��x
G}�nrb������D6�o-��t����j~�2iL�$�!h�f�D�cXi���S����,�Ӊ�t��^n��Z��=Y���\�<��Ȏ�*����x!�:�z_x��X�	�_f��N��+�=҅�Y�
�w�y�p���]6U�:��){҈8l��G�?��9�K�� f$#? �V�h�x��r�Y[n� ̽�m�5`=�X� U�]��=y�+��wZ{���rc�ɰf�ꢖ�:֍fFy�b��#2O̽	�\&v.��LɈ(O��A�A��Q �;:����9֕�o�pTԤA�֧x���V@Y������=��^х�ɀ�Q�B����ՁƳ	�		�y-��}��Q2�sg43�d���z|�׷�Ia���ν_��@��3x��ȫ�ˬ\�ܽ*(hB�ͭ�����6�`uX��r���p�m�Mn;%����7����oM���{�s�a��s,,��5А�!)Wq[�Pw�l�#��<4�f�4���&^�R<���k�v���&�)�ĎY_��/�U?��K�S�>7C��JʅZk��Hn�=`�L�m����'tm� �/9�B�?F�p5s�7=�P��:�R�tZk
��e���� ?������M�7Iv�GA�cu��Y-��s\é�aJ�س��#v�)�����4�w�J��@�`�C	Ry���{[m����S�$��*�/�Y{'~����p��4
SE}|l<u�4s���<�-��/��;6�̖}�Du*���J{.�TccEP�-J	es-}N�w�P�#\c=��0e�f����]iXG�.��2���';�ֽ���NS?epaդ�t�u�����=�%��J/��ɍn��zh�Á*���� $�ڈ.�����!��$�*�<�N/�[� 7`�|'+�属���9�ЄN5z��;��||� 9�'�W~��]ʣ!+�ݙ&Þ�:��AɄ�K͑����p�O�׫�-����G���D�La؟�JcV�]�%vM?g)�9.:�ȍٰ��I�,����OS�e*�FNu�d��`��T��/`x��PT2� �O/��p�\L�Y�J�Ӄ��Ƈ^#�����g�l#���AT�����3Va�|�h�-{/�s���,�Y�rg���n*Q�|L�=]9{��T�IT��b#29�����6���)�-:��@b�x���H:ڰxU�Q��p�1ڻ�N���ƍ�#h�Zw7{x����&:ϒ�k'N4�m�Z�q�/��B�WQ�H^}�I�xP���N �R�c;�ir��hjy ��ʫsz?5o#ť��b�l�!=�")ͣ~J���^E� ��>6�7�������q�h�9H�� �0���������*+��e!]}t5_
Ţ{���"} /���4/9�f�idBtaO{">q�d��KoĒ����ܭ�a���P%�{o�k���> �.��v�#}�6�ⴿ�d^F�;s������=m]R��:�� �-��v�D���S�I�Jp8Lz�ɠ�K�I�P&p�pVQ
5H��tÌ����y�$���ZW� �ބSܙ&�0l?'���l\��
�ꝍ؉|t�D��_>����ݫSB]������`��k�7���`-���!�xo��6i����Z��#HߙT�4��͝=���am�����P�����j��U���`L~?���U�}4-J[#��S^�e
[�YF4sq�Hde��/��qW�?9���V�Fq��&y��o6�ʓ�%]#����3H��z����f���a���9x���f��E��:_�=�|X���os�U:�!�Dl�]_q�+�ӻ������$�Ro 8T:������.���eS;�HuB��qR�|ߕ�,��g�X*!��&EW	�ɆS�L)�oN��W�K��jB#�ͼݾߔDGo�^�y�8��Q�V�	��0~����r�����hA��>��������c(lz�����# �����T�5d	7Vk
�Tt�$�;䙃�� �?ʥ;��4�v5>A!��|>a�>��<2�4:4��u�MG�z����=���)�b�� Hy4��{n����P`w�a���E��D��u���{CS�1 ^�� ���I��!�A�Is5%��P����r��w�.߁�2#<����[p�ހ��S�L�hd��-����%�#ߜ�2�3��)7��?��:j���3�y���=Hǁ6��K���,n�n��p=Q��i\@�A� ]�k7��S�;����ۓ�����̘���ڒ��6w�|!3�����@����>��n���#O��'[5����7��rS�P��Mc���ELeB���P�&^��o1�c~��n�,��\}�z�_j��$�0z|�Z��J�Di�\��N�}�[���\
��=�gw�ZR�h���q�+�7�p�Jp��P��_i1�pl%Uh2���O�j����=|�}[�r$�.׀醭�Qn�����}�N����>�/��4K��´��}�&C �)H�!���Q+��4R�Ǳ�c~a�J�!*}&��h�m�c��=�xC@����`���k�9�V��V���IL<��������J��7��r�}����ò{�5���N4�M^��Vpi�Z�԰:9Y�9�_Z^�t}U�oH|(������
k3��?2E�k���k��s'�5#��uPL��G��\��&�M�)���ԧ�YSH�$�+¨V��7�]��}�J/j���G��ij�2!F�$q ���/�|d�}p�!3ߤ��5y���|���%�R�vNt{�i���l�Z���J��ᒜ����B/,#��ʂ����O)��ڋ��,���y"�c�N��z���Ґ!��ng�}��";�;��+:m����a���%�,�*-���#p�*	aFq��M����*!}��ߴ�/��x�]��@�N�^b4�v�)x�����8�2���(1�5�ǜ�#��=��K֠��av������I׃h���>����?t`*�ddҙ>\<����4r�g ��)�G7y�5z�*��Aˣ�\�_���5gҞ���ܿ5��H���P��Ӏ�M��K��n�碇	娕���L[�0A�K���	T�g�YU���i��\F��ɼ�j-�R&u��:h�`���F��eK)銒�j�Z���z���2X�	RY�T��7� 3~�d����v�zKh}n��A���6�ȏJmK�� F�`X��^}N��|<<�}@���D�˚�| b��c�a,_רFl���Y;���"��O�u#y}]~.J*w,���'���X��iG���fw��~M3%<����>P�m!�:�U�n`��	qx���k��)-f�Y���y�5���.,4�!ﹸ���ev_,H^p����0�Y�3��)����a�O�3��K{ܽ��o�#�(�����������u� =���&��0\�K�|�J��\] %Q�v�+Q@���i���C��O�\�6���z��>�˽�`sjqK�$ʁ^�x�A�_R6�c����'(�&����jmf���͘�p���h��DW#�#�ɤ� �2��L�{C����w7����Θ��~N3��b�$_&ODG ��!aa�L2�״��s^Va�MAOS�� �У��K���Y�|����ɭ��� 6Ӡ̨�+������U���9>
�[��tE�s�����9��[&��מE�
S�񈪭_����A(4a��eG���)��a]o8�\�k�Ow��g}��5i�c~�����Z�pȢp]K�J� Mx �`Ů��,�Sj��2�� ��vk����Z�|�f�O��5�9����#JM�)�o���TX��u:6��Ϲ��#���8H��=^9���,��xmyɥe66�������Z%ٯSb�����]�M7BE�=�Hf�Y9�L��/�P�pq=2�����f���L���C9��~y�Dxxf��|[��8�6��������Y),�8�ܯ^v�&X�����w$�G�������F���P1\3ҥ��HC�Ngc��J�QA�h���](�߫X�zUy�l��3������:<���s6��<g���#2��<w�q��"����|�����!:�#�4Yd��:���ڒ U��z��3p�������/6�јn)+�](C	ޜEV��:�a'���T�H��j3 ��u��BE9-�M�h\��j������&m`�y���<]n>���r\�.tg��\�;�4����X)���ڂ����X�Ζ���)���-}yG��g*��8��v���I�x�ƞdܷ�HN$ZH�R@�և\8 }.�s���s�Lt�7��3a�/'6��DRlz�@�z&�ѝ��Z@9�!H���
Ry�)S-�z��oa y:J�7��@�,�C&a�Ě�����D���V_�;_���;9��׹q<��+���/Z�����A�PH�h}�M�����v٪��b*���E_O����#-݅z����$�}�����q��{�Jej+��87l
��
�b�7}��]��O�c�g;m���-4�����4k�H�4,2�a��Q�j�`�rP��r�Ιd���1"�OJ����Q�t���u�y\����O-H�[���Ӿ�Q�;j#�✓������9#$���[<�x�s�����8Q����Np�m�~z%�냣��y&O��	6��p��[h+lzV�A��K��܋/�u;�c,��g�9���{K7Z\�"�#�ݘ2nf	�����-�֊u�h^pV�,����o�Xr§�Q�Ѓ@s�E� ^~�x�ϕ������� �9�w�@�#X���{�����)�-�l9��zf�(��L��ˬ�UI���D�{���I��PG�6�B���IQZl�a�F���袺]C���%�����,�G�AL��3Dm��Hw�cܛ]"�ɇ7
%��L�W"�.�� f;�N��N�|��K4���L#��	
�3 �:7�;�X��9I��=�A<����zsX�OBsB�#�$ä������,_cJ�b��Pr�d���4�}(h�J�1�����%`�'���<��i���P)=Y҈+���Z!��m��UM7Q���E�]3DQ��n�����fU�Т��s��n2�?���z�7C�Mq9:͂z}ڹE���ׁI.���~҈�t�P�sH0�ZQ9����Շ������[�4eHhB(�%6U���=���|�`���a^��:}L�W�`�10]�|A�Dj.#��x�����q�zy��}s&�,�g�c�)�Ajo�$ ����Mi(+0�Ә��c(�� �qr�eQo���*IJ R !XsْU�cM{|F��}�R�-PŒ��@R����ʄ��-ڕy6�'���Im���[�G��m/(��A\����I�~~�:��߁E�!���J��#T� i��G�<
�����J��㝖�����Wmd&��H.ع���ד60i���'P/<̬�� Q�=u[�{x�7�/��^@,vo�ϡ�s�4?J�D������/*'Qӻ��.X_��ہC�I&��j�:�:E�jE ��h��gҜӒ=P��Rӏ�o]�bH����/Z�/5�o�:F.~�!�����U� �X�v4�f���Ō<��6�*�ZJr��/��)&���h��hE	����"���S4$}�EV)��B'��-�R���2?f4����C>�~��`7fF��km[xD[Y��$Q������0��Y�:��ab�ʹV�u8X-�`�DN��H�P���b����m��}��M�Z�}���Ƣ��ÓD�	��ֆ��\�\73wm� <qA���kmuպ��/�u(QGO[%�ߧ�$��eՄ�g�U�6�B�Vˉ}ii�𤐡��⨿������_���n-|-��>� ��ge8�T��,�Cvqo�m \d�an$+k�X0҅�=�EK�[��x�4��)�&Z��?z#�'}0+L`TVټ���j�`8���$�x/����L�,�ƾ,�X$��3K�I�N��VWQ�����Ƒh`ev����#b{L��g�ecyT��ֳ|����(��B{�=q�f�Zg��y�����3��Y4r��;G2uQ�����m�;�{���#zt(O�����S/ds�E ɰ=�(c~�m
����*�+{%�΀
���o�~�mbg���Ͼ'F��/;�P�=�V"A�%�m�i�I`�*B��Θ}S�D��5��9���Q��C����I�1֬k�����1ܖ�s�q��
�B3y���%�u;m>38�~ID�arj�5��/��5c��'.�-!b(y<$�k�1���[m���K��t;;�#F�^ga/�4�;����d�2Kl(a�9�USi���[���xM�lT6a�3��8���'5��7S|�M�S��ۆ����܉.*�f�'���9c�c|"ߧz��{S|�<�4��6�"2�@�
�r����Ah��߀�$�!�Jq}�F�*R��7d����|;i�m����,u��\���y����D%9Ϡ�.Qַ��L��&��Ŏs,[������X���Hq�洐�¨K<U�z؍ȶhBKy�rP����n���(g���.�tG~X�qbJ�Q�T'1���6�W�}���(�@���Yh=�
����ď$���t�m��T@̃*-�he�ss��<��0��N�duSX���+���
�c��˵�`ٗ%��
���'f�z���B�A��@%/��	u|��Bl�.E�W��ŧ���Ҵ:]��,:ؔ�Y���, �J�@�����ҝ)˚��Y�
@�+�@��ˠ통������K|S��\: Cҫ%�硛%����T�2Pw=4�4��P?E��;�qT�z��	�;nO�ċ��N�{����}tr3脃�ͧ�pr�Z!�aB<?ǚ�t�Fl�G,#.7��%*���N���u���S8��V�*j!O�GX�+]؀@�}:+E�c�7ǋ�@Qi��)Ψ�G��~�KH�� C�m�F�)��yb�R"����ㅽ^@�y�b����D<�ɦ�U��b#/����+��;D �����ׂi@���,Ee�vl�W�r��W\7	��%����i����d�&/�Ȇz�}Hq����Y��-ʬ6���{})������r-���K�k�.6�2��6z�r֕����,z�R����w=�/� �zD6�q����K���m%���ɢ.@�.�����[�Ȱ����s����U����:�2��z�	s9 ���l��I��oV���:0���j�����]t��*��qb�'Z43�څR|����]�>����AjI[qW���u9����SͲ���v�	.�5'mfq���ȓi�!�pݷc_�~!E�}��DS���`�8��Z�p)�*imR=�d���yo{�F��J8����S#tF*����P&qM�^���N��`�D��œ|�Ua���A��S�j���*��4Vr�����_�}�Iz��ؐ8(���*�%����%��ݠ��ٚ�w��z_t���@{2�4=�p�g��Vd�JdZg�
t��)�d_g{{��U47˾;0� Ɲ�3:5h�w�$��gY�@9dz�W8��KQ�:P�x����-פX:R���J8{�cb^55��~;��A��=�\@9}m���ۭ)���\��}�@����[���	��R�Z]eeL �[�
"����s�O޼&k��JB�,�VꚚ)�`Q%�a>��;S,��f�M-�-N��i�Ȱ�-@��|�<${k��RC$t2[07�6���>nS=vv�
>��̣t�T����Q�G�Ў}�[f���c�v}��I/���:�)� ��oȻ.��v�k`�!��1ؔ�5
�L]$�_��Vap�o�z��3x�h�FGle�YQ~�~�O�����h@�=�݋Y��qȨ�JV��k�V�׮�L�U�L �M��n�2P7��љf5_��Uݹ�RK�U��V�t}����V���"i#�����u2�if(���qr�0	��D�<��`;|7���oN�f�����ގ�{z�2��,�Cky�.�Y��MZ
��s��Ul�֗��]u9��\7姵ɏ�>ZN�de񪄻�;O��K�M�C���@����j��o��,N���M�o~��^�%��D���$�����6����:/��η񨞰����dۺ܊�,VטH��Z���D��>�_�m��b�	 �(��;&���
�zYⰣ�ih �����?�ϓ�#PR!�_ &���	]�R�C��W�Ud+ �24҆�-*z��X���s�qaN��I�wm���7]����Kh���PS-m���7�Q�#��m�CY�z��b�~1c���L�]�zl��G�,Y��p��ם���
��o�8�|�-��'�@�#�;��x���A�يYo �j�4|`-#������o�oŝ��R*�36�zю�����_m0�]2{�-��.펳\�+oW��h�}�f�>F<.	w�!�K�����E�\|����7IV��+�������݌EQ��O��՝�ր]�<�Rݒ )����N��^����{o�6r�����T8�g$=��@��g;�Xr��I&�h��� ψ7��7��g��9{�#O�I�!1�n��Έ���y>7?1�%6z�Dk��h��E'Л[߃7^��7B
cz�^����ě;7;#��h��a��߆R�0����t�,�:��6�4'���oB�y*K��c�����x��s�zÉN�G|��v��|B�a�g�PP�bj��b�8�7���c8�"/��&�@��X[�k�ݵf�;��sm�*�9�3B��mA�LB2��MqN��#?:H�����K�2��)�ͽ��g�Ǵ=Ww��&��ӿ7l�ʂmy�LPd1����3����{􇴷�L�����hA{`���"�߉�1 
���U��}��1Mu�(�NX%"��sm۾K����~f�t�3 ��()x��xg�h�����:��p���7�����Z�_�#���}��X����40�U�Նv���SP&���J���$��<�������n�_�%�y�UF�ѣn���@nɞw�HP��}n�H�Y�~�NJۣ�)c�?[k�X�h;���XA~0	�n��[!�����q�`���/�M �4!��7���׍�FRc�z��h����k?@�r0���e����l�V6u�rl��K��W!�g���{�#���D��ť4���H�q�ճh��%r�y9�b�s�Ӆ_=K��� ��ڻ��x�*�sӾn����S�Lm�u���g��!gF��6�_}!��5CYxI	ҙ\x��5soٰ�+�]Ns Sx��(����+)�'O.�քb��Uτ"��[��Y ��aH���H�C3��Y�.C���C������P���e��qw]1'-�xg�ʊ�_����t�x��{�F?X$���Po��t'��dAk�kl��� >��P�V-�?ܡ�?�|2�5��6��TA��kË{��_�A�n6?��'�j��c�F�(�11�8���K>;��'n��U�Ev9�eb�i�b�����2��e�8p����G֩x����Q�H?p�N�D��wj`�ƩP�'����ϊ�7�MNV-�F��"T�[�W#���s��=*�?%ow�M��0V��^?���E!A륣�?D��<"���$�V�ő*��-\V��(�~�N8pq�&=��r�7?v�k�6J-� ���0�K�C�ϓҕ7�z���-x���yd� 5���J� �>f�I���V�Xy��?��K8��(�V�F�	Ր�DU57&Ag��K��@���������;��3�t(�������|��4���VL�a���7�v�g���lQ�ѥ\��^���q���2�8���Bl��#��L�C����i@Q���Џ��솞=�����W�:�gd:�rJ�ѡ�.�nP�Q��c��T�LO�NK��*0-2�Gc��g
�\F�F>K M�����Y�PZ��\�m�/�`��>�Z9��#��8���x�iP�rɀ�4$.���rV��{�ѭ�&�g��]�^���n�wq�xO�x$h�Mf�c���L��k�#V��6��\�[�<:t�ND�c��*�2N�?����wBE��MaW@c��:(�Rp-#���ȜM<J`�剨K�CI���H�¸�/���=� �`I��䉠�;)��k��m�.j��G-�3:���U��"-�Ʋ��m�Җw�H����q�-���DpS���
-z�ǖ�p�ܑ�ԏ��-ѧ*-�y_�.נp��Ju���q���4t�6-V�����"o��C��I8>��>2 S��R_���C�Ɣ4�\}q*�I���BN�d0r'DwX7���|Bg��F�� zs�h�V�Ω�O�O#}�����͟���BQ��g=�����7ey������k����
���ls۩r'����ʂ����o�����EI9����Q�jxE
��%�;E�\����ߏ�q��g'�)B�Ժ��VdI3�4���R�\a>�I7��w%�O$p�%	�;�uMp�'����C!�/4 ^g���}���c�o��Jf?]� �J�~sw�N��ڮ�'��A:S#3W�c�D��uQR'�۬��3�VG[Rr�\���ǥ�4(s��^�D�x�-W��ď1���֠U�i�y��e��,��?ɓ�q����Q��]X�nC�@����l���hH��R+~v�P��
�e=��{��	�����5&�_����J$:`����ɋ�N�b,gt���7s}��/9�$��w�ȅ336߯|�I�uTJXD�F��yZ��>�PG��{ye�y�v��q�7\O"ڐ��(p�̐��͙X��ʂ¡B��<����r���
8[8��V�A� @���p<$�-��5-�Q0���4��L���e(G�Hi���Ew4�t~Q���K΅e�;m]q�t�G�0��B�D�E!�,��b��n�X@4��kI��Q���6 R���t/1N+_6k"B�&�����w&�)d����;%r�2t�g����g�ٹ�T�Ё�d6�qr�Qzm��m�5��&�<}�}��a�deQ"�=꿆�4���1e�7~�"`gO��BN�a0�\IDo��g������	"_)�#��8Ǒ_�W���)�K���;C�z����VH�?�Ocp�e���nD$p
�'?~`T��0|V����0�r{��N���d\;H�����j���!G��� ��N�S\����:P��Z(�x�QݳHp���!�C[S�fq�>�S1���ag���6��2eo�rŝf�\F�T�fֿκJ�|��tL�vU9�����"�V�i�����ύ�`p���Kr�`�� ��w��JTHN}7J��5z�k�k��<&�"�N�����7�ͭ�:��j�v(V���q~�K{�'g0ґ������K�8�!z�\�������Eg���'�-[���>0t����G��������}4_g�ʎf�����$����G�(�	C�G�st�!����c��k�*�E�E�������aż�	J�	�ayZݳ�M1tc��t��E*�m�5��No���8��$1����!�J�:��X�x$�д�v���r'j�C p��]�#\���-��b��gMDn����"�Yp�(N2�n���� �37�-��ٓmY��S�W]��U/ao��e���ŏ��C�t���8�~ڈ�-^��H/��<UQ�v!�͢wم����I�{��	z{�If-� ��*������D� �4Fd����pWo����v)��n �搷)I	��w'iv���%7~!���<K�qW�J7ۭ��)��F�p���
s�c��nnFk�/݈R�On���q�2�w�I
��;�7+����+*q�>��O������_�a7c]~5p��HGW�ʽ���4��7�Y��z{�n�O��I������?[����ћ�U3K�֢u�3�}|���%���,�"��쓻��3eit^q�L�h���؜&�=/��yn��%�hr����zO��"�{�v\-e���iN�B1�	�	�8�l�����y����Ub��҂m��b$�����`��c ǣgwb�zq,u[^�gQ��\	��L�f��	O�%���ѿx��-��gߋ~"��$��
p��z7Ѡ��<X�N�=�TӃ-H�(�g�1�t�/*�9���!"��^,��"�a���zU�:�����~/���ةR4������&SpL��z	��[s�G ��ڝqO��,T���� GwHR�9����&�d^R�[�r�㮻�u�o��q)z擇 �����Nq�p�+PmRf������\�����sՕ�[+[��L����n�%r�Z��?�ܦ˵ַ��-�wq��t�><�p����}�٪У�g�{����F�� �����n�/h�u�﫹�-Ķ����D�>��sC?R�y)_�>~�㍰O71Aj�D�O[��;���x���Z�22� �}!`�7�ypǢM�w���w~ T��8�����\ԎO��I�����Ix����MkU�C	Y���a�֠M!&φ�>E� K��f�����;��[�gJ9�o���~��/�솨Ki'm �HUGA�[�*�ܴ�觜ЏA�	p���E��u�i�`�Sܘ/H��A#t�89�<������ll?�1�U��Z]셪2�����VIs�de�����~ꙅ-�����G��9��{6�r�����qX���6ԥ�p������+�<�Y:1��d��H8r;�f����!|�1­-Ek2�W�r5>�Ęε6 O��dJ6�s��R�sԶ����B����N�.4CO���bi�:��9����ɛf���O}P������\�I��H��h O���k,���;�5��� �Y/G1�d����Pd�/�V�)������2�.�n��K����n�Z^�FJ����*Ւ�7�	�����9y_�B�o�o+�s3�kӖ��
Z�7�5�Zv���7+p%$�Hm9=�A��ZN2W���X��1��A���z
��nߗ�~��ß�t����-�z�~C��l̥�fEڰ�*$���t�j��? �p�߻l���0�V�1�(�С�u�o���k%���rp�c����'Z&�R{N�h�����SF����n�vk5Q���)�|\#��$@�n�ANև�bc��1�βl�ֆjxA0gE��U�o3A�~W/�8�b�!��V���	�P�`��~�M���%�$�E�&:��#�>�T��K\�������В���Z��&ۇv����%f��f���qx�n6��n��
�cl�MT�;�(�ݟ���E�J��#�Nq
be ���ߖi���~���L	,���E��8Jz0���:�:��wo%L�$ͯ/��,|� �;��T�W�E@�wr��]���9C�i=%�ў���L"<~R��ѝ�	@��	r��pai��̡����p`���a���F�*$6B�
���2s)۝��-?wi��M:�4�ѣ�w|!�xf`���f׳�4������̢3�
� Q��f�-+[H&�%����g0?g.�ٷ5�~'7`���"��r��ai��Z6 ]���ە�������V�����V,�	)�z��X���c��S�1�!MS:��4�C�.�C���Ht@��>M�&51]@y��oa���(�[��"���H�(����^�[��7�
����Jᇨ�Y1�F�2TlV�r��C|�CW&�&�a�?�ϖ�~ئ�Z1πU�N�WF�*��r\c��OT�{���Ra�����^�
P�t��/�^iLdn3��[��>6��81�=n��[H��u��#Y��ʆc��o���HE��W�̣�)?@7~ �-�>��4����E��̀�On5։͸#6�Th�+��7:1vM�,U�q|2���LD� ��v�X5J�ku�:��]��$����ws�HE�l3%�O&m;����p_[�fr/w�l^����i������"�n��88�'뤗,r��Lox�N�ڍ(�\�Q��,�c�-�1P�����Tشx��u�K����0J����z�3(f�d&�j��0�F�jR�F�1Ċq�i�����(D�;��z
��YM�]Yp���8�:k���"UP�>���%/�_R�Lĺ]���k�x��.v�;��u6��de`�)��}BxЁ���;���'�N��|0K�O�㏣�%G�2س+~���٥�E���VN���	�9���l�]�<��`�G�g�4ȝ���#��TŌ�2��z�
�O\�Ҏ�IJݩ`U�ؤu�WF%�v{/q-:�����]�����Vo��Bqk���V5�u��4dgȤ7
��$�{�r�B|�����\v�v����ղ?�9N���J�P�%�1I��E_Ո�	��Th4o|���<?�2�%;@uq&�P���[��1�'�v�S�H���n[v��a�U�JZ1�T�ئ����!|�����:��������U��X��A}b�ҍ�ܘ�J�a�� h�hA����'r��d�K.�0J�s[�!la�q2b���O�����a���/�ږ �� 9Ƃ��0Q��:b�g��F��t�PM��|o�W�3aZH�d�1OK�uh��o�:0.�����MN>]�?u��z[km05��JK�/N?�(6��H�����~�V�{�f+��r=�F�͒�3��3�Y�j�+i�;�i�<��� �1�w>Ee�pp������_�ܘc�?��8)!N���5���XHaa���Q)ux.�<c��Y��Y{&�RZp��q��`�Y.�Xm��H~Q��sg/�7��B�+m��ؐ�o�?����m���`ױ0K��.����]�r���؄K�8��e��f����6�vz�oQaI%���r��"��!O��6�
xH����S���"�(���c��e��hi1E=G/�-K��(5`�����0%�������g�_`;�K���~�u�X�v�jb�oyN��m�lq/7�acUaF���6��q��ʘ��#��z��������7�p�&����S\}�T�$Ռ49�}Ʌ���Ư�F$h(*�*���5x�z�[!�B���_���uy��(���"�)Jו�R7��a���Zk j6��GG�ȣ�kn��9��)q̟w�(կ́ɝ\=2�M�](3BHe�`�tc}�i��Lɞ�� 8ED���?�<��Zv,\�#T������t��w>\C�w=l�;�WV�P�IK'�����{
c|�Y��+X��^���x���js
2�	��0�)��>�d�i�I��:��MD��T�ŝ�D��,;�;��]�m��I�B�B��}�4�l��!(@��}�b�q2n7���+z��-���fcU��dK�7hO
�U���;��x��F������=�L��X�rm4� �a��M@s��O�54M" �K1A�Ho�<����'@�):-�j7���a5��Q�*��;q2JK��67�b���r��І��!���̷��hT�uC�DD�L�����H�u�SVs`�*W���̯�'w�҅��� ��nr�嬴{E�m�&�[��T��5a�MJ�䚨�"l�`٫46��O]���I�XRU��v%ϻk��������	����� ���#b�H� ������B�>9�$�-���V���C�X������@,�A�v�L�3| ��*0{�q��-����M�oTF����:#^&�|��B��(p��uz�_���o+���"�~���x�;4^�=Q��pl��y�};7@U�5dÊ��dב�T+%1ħ��4u�x3���.D�Uua|Qż�]�y�vÁ�ӳ6Wo�k�[^�\M����y.��xo��?-�#.e�� �I�P�<p�vŽ%��a��+G>c��!���߇/�;�Ì>}o��b����|�w���[pt_Ma��ꦎYWh�$U�7�$~�ҿk+V�1�T��K�?�Y���P�^ƃ��4$�5��]_�f:`�I�F]�O�41u ��ߡ�-us�L~Y�8vi�%��~독LxT�Ӏa@$�>��-�õ�C�]#^	D�^D���4A�@�WDG��� !��ohHϕ��:Ҁ�Whd��Zu�"��29<�	���0F7��If6I�h0r�=���މrɰ�9rD,��l$?�C�$!��SQ�����	,��Z���g�AA�] ~����E���X3�g5 �����:I����Zd���8B�N�!Rl�r�T%�A�IP�����!��k�6���[�A�Q���V�p��')V�-�8N�qA�8�g�`�����Rgig�e����cY?�U
��
or;W۸����f����*�jѳ}7�(,x��uw�W�5j4]��u�9J����4��R<	�Hx�)5HS�hF�}�Ƽ�2�P��dM_F���7!&{�P�'�5xlh�jЋ����Ǒ�Q��W�-:�3%�W���B�=����_������ԡ�hj^@	��ߙg��/� �=�;�Y���$�������������t�K{:	��AZs=p]�`��T�Mɺ�	��Ʈ�4	�1!�<�Y~u)X���-=o�:��X)i3@[�����:��D�m\���>�6�����_���p�cp*�k �G�5K:�宾z��΢.��5(���E|��j��Q�m�O=����ӎ�>gYo���}9���ʃG$L��C��F#$*y�z����}��^V����ϭ&F��G���6$� 8�t���h�@��}��M���۶_�8�9~���F��뵻����� (H�CBX�6��6r�dq�G�#����D��V��..E�5΅��FD�8��
-�,�]�����DwoH'd@7s�,*;@��fJ���t��%�J��\!�����.��O����5��EK����:���\�^��!�}RR�윖y�@��W>�mU��qX��!ޜ5-�)��<����j��� �i���}׋"o��Jdx��GX3X�.򛙐�6@�J/%�3�vzm�����J'�1�[��ꘝ��$��2��ㇿ��W�w��ۜuۘ} ��� ��<v���-��4���P�>�v����lp|������c�?���D��i)�5��Ի泃�&��+Ź�*!������Fg6�N��q�����h*�X"��]�x���x�����N*x]���Ȼ2�(���O���E�9���Nt�O>|Yh ;��M�I���B�R���d��"ǩÔ���)%�����K��I ��������~ܥ΋8y�nV�8h�k��WaJB�3F����C�W�^��_�@���M�}h@�D,x�+��. G�:���ǽR(��ƼGٰ3K�͡�sV|:����n��Ö���Of}���y}\
�a�;�����w(�пe�y`Z�-�_���1]P*��-�:|�"����G�����BuL!ǊW"Fc����봏�zY�rɌ �g7��"�*�㇊�>��nhuV�*�`|�h~��s�<�$����c�v�/dX��T�f(=�7�wt��}@.�4��ү�+��]�bwl���Y��^|���ް�74�m�E;�Wo�wR�u�S«H��d�}�.�r#�����,�,O7F9-���%қB)3��鷪Z��LN�]M�ue��pG;�'��w���n��T*$�pb�_Qo<A�$�`�����o�;�Ï@Y>����K�$/�$o��Ԑ8��
`A��"f�;��Ws�b\������y��Fb�@�$��ֿMBr+<�kb����*WI�a�S� ����+��r��'�W	�޶�ͷ+����ځ���a��o̒���f�V<ΝFU�=<��iz�F��pㇽ��8ڄίl��rH�aK�t�'�䛰�&2I���RK�!X���1qE�m�W�)`�h�	����y�b���0��vG�{����Du� }J6�m���aAi2r��FJY��sv��G�oJ�}�N���nU�S�����N�@���[�� K@O����hS��y��)	�:`�fM����@�d)��q�W��3�y�3N���h	�O3A����o[rGz�{)����C�V�Y����D�P|�>���/\C�8�'}������D�M/���QЫ���]�m���O��}�v���d��ݹ�B��C�<}��@ ��9�h)iϥ�V&��d������x ��Uä���.E������A�������ka�܁G5���O�h:{���&��\�63=��]�WӨW;��\4{���:�(=����J�W�R܏a/e%;B��u����`�Yqb����=��<����<����Fnxi���(����Yyj�"�丑�V9N�Lݢm��%Ր ۸�wF�b80�כ8(lr����>�i�c2geֱp��U@�ÃPG�CL�����'+΍��#ކ��J|W�8�kx��<Dm@�w�Z���N�t2.Kt=����/�4�"�b�)�xQ�n'K�BF)w�-!W�Ł�����r	jK�VI���=���z�QR��Փ��0���xG��M^*?�,����� H��h����^s��.~�*N~-H����ā�1<pk������^`(!��O�d�]���~�P����h�P�������. ��3�WT�= �%�9^���-{(JI�T��J����\��#�R�8�0c��,#{r���{�a����y�٘�
��n*j����I|��'ZQ��K�� �a^�^��ί�zY�W6k�����p�g5��۲Umr�:����9������b�&:��s����5���&�8�Fe����!ȫ�^Y}JFKF��"�
O�$�W��%{!E�x#Ԧ^���(*�����̣�D������mӣϏI�\���m�԰�h�˔���0<]�J��2��{�t�(�^ܤ�xx�S�)�;f)Һ��H��$L!�1c�p�@튑4t-����k���B�'�ׇ�JP��r� cU��}Q\%Ưp�=�����-�K�;��m2w�|m�bI�)����]nI�j<k(J���a�X����A9A#���D�>*d��z��7Z�uԇKC�	��߁���j�$�Էg-F	%�`?8=NP`�74�%W��S�Ⱦ�f�_!8�9Q��j�ʃEC??�j/�0���
3Y�n;X�����HPD��K;`9�L$�Ψ"�E&h����B�J`	{͟ѫ.y�r%;�t�=��9���z#U�E��󿦴�q�?,�"�e����	R��:�yY��7�疦�Ԩ���?~/�!;�?�crFN}V�� �)�Bg@n#X��`n��aj��x�֦��/�x�>��#M/�,���ڱ�tf*{-1.�Td�߉δ�mj1�q�mU٧��k�-xN�_o�5�C4�Ae��fZ���|O}Ư����A��S�0t��f����r�"e����5eB����)}k�8):,s҄�[)w-������qǩ@%"�l{C>k���w��Q	m��P��0����ރ��lp��;�oT����IΑ���ﴼD��,����'�dɇn�����Y��DO��;� �Yk��C}���p����#uu�i�a�F�Yw�!�'ZD���G��R���!u��0���Vǭ��[���F{l�r;�L�����3+�x_��[�v�d�Rġ�5��h�.a�y� ��ȓ8I���`%Ua���'��4��n�dz�z�o(cKxk
�E����7��N�D�0=�4�M6�o���4Li�Q�Z���CV+��S�T_�����	�b>J珢Zk�ch�K�晬��݋����RF{�n�wČʾ3Z�w����ҥ��B��0N��fq��mr�q����ذ�'�ݬ���g�`�>d�c�#��/(��a���jKU����ƃ�)��9��mg�L�/�z ���X"��?����ӆ~�Sl�vp�'#�Ea�dO�l��3%C����	`�V ����_�w��n�sJ���K�2�#�K����E� ��6���p�o��W}l\���k}�_�R��W�����fX/r|�%��Y��	�w�oߏݯj1%��	�M�<�n�?�r���/!<�� ݫ�
\+'�kb"�N/�i;[HM�T+��/3S*������+*�31��+g���5Y���ȫ���b��p1��I�@ps�3v���N\�O�{��\�����O� ���3�*��(�1p݂��'+�?!��qF�:���g���KAj�)&A��7��L!*E�y=hE�W�\_��\H/HOuw���q-��r�ne��}@_���HoS#�z�g�Ǽ��0Y�m[N��U�H{�������:���Ф����jÐ�o>&a3��#T�ؘ�t:��8,�bT�j�3B�yD;{8�Z^I�\
�
�>,��ޣ�[�i�÷N���Yk��H1��B1�B��M)�e���+�[nRꮴ�d�PD�|vR�,�������TiW8�n;��7���`�G�tP��%�������ch2��'��#��U� ��:;j�IE>��)�.�+���Q�`?^g�6�*�X�!$�Q{Q`�P��w�㜯��Q�o��1��E��gJՄ^TC`.�o�C��j�hv$���s4��_p+x$h[���D�,�Pq;��[�k��I�&�H%�A�#mOV܈���=����V�zGr�SF��JE^C�=5#I����p�߬h�DxҪ|�=��&Е@�c��Hx�j����{嗗�h�a"{��e�c��o��T�|h�]��8��a~-2�f1F\.-zn)���_b�k�xq� �����δi�Jw7*q	Eر�
���^�񨧼�H4��`�A|��^<lrΚ7�|�5�$��L�9\��5����@����+��#d���h�
������4��}�Ǜ�
E�@�|�G�4>"z	�T'��ۥ�0c�"���1�s��afnY^�Az�aT�k��\������
��t�	�`R��Ic�����sM�ʒ���x�/��_&+��n��8f�c�<���,n��-����C�@�犂9z�%0!�R����3���ٌ:9��h���@l����>u�6�Ĉ,aB�|�W�ʸ�����_�֣����q��f��
Ћ[F � T��_*���0dlS���4�#K�lʹaL�Jsǯ��H��`�᪰���P��.����u�P�]�{y�֠O�/���_/xf��E�S�eS�&����\n����2�0��ll���R�7_Y-s�'�W�}i����9M@8��	)���}j�]I0�a��6Z]G"[�P������&42s4��b�w�1�R;�H��:Q�Wzu\�\�qID��+��с�L�-y���2�!�Mb�8�4J(l��<��Ȑ ����Z2���n7�Ȭ��'z���$J2���z��`�j(�I/l=KYB2<W�Xz�@hjF����SIy�'��vg�J��ٲ� �&�h@�-�L���]�o��͔����S�Э�(�ْ'��O�?�IWjơ������Q��T���&� ��Ĵ��I�L�Ȧװ�����ѻ	�2�v��ے�ϸA����=
VH�̀)Q�V7�x@?
TK��������7�H���ҽ��U���S	����X��G�֩բ��<NT�X0���cr�z*�9�`��$XZ{��ܓBּ�� ��#�zf���}TXe ����Q$U<[<�nY�}�����U�������wD�?��Ii�OX>�qIӪױ�0Y��ϢK������1	�.h�U�7Q�a��I�f)��(RδfG��o�}��:y�&{8��D��z6�2�a'���@�L�k�)�{ꪝ��
�<W�4�q���
6|��.���Y��:�����$�xkEy�E�{� aB���F��c~��#�ǳ��c�g1D��k����T�Y@�m{o����C��,QҔ�9n7䅔h��u��X��W��w��|ȳR����
l<O��A
��5�'5r��{�Ynd�,U���A]��и�דbY9P��~q!�&���,�+=3�K?����_oT����*u~�p�� ��LW؃��t�Bf~W39<�cX[����q��F3���S�\ը��$�>:�B��"@�:%�sLJ\c��t�!L���7z3�x&WL܇gw���;�Kq�e2�$M�Qd�b���^m<�6N>f��i��1���V�R+�Le��>�.����[VE�rs.jaȬ!L�u��-,"�b�H^x P��*����V[<���[�4��m!��hQ��G���ڛ+w[V�K���x��FL@�س1��7rl���A���Eas���!���~��h0,���r��=�����$��'�hm0!T�
���<���*7�;�@۬V=|O����U�fK��	4,��S��T^�U�^e`a�CVZ�_;h+7�5*�Bz2��i�-��@�79�����5_�8������pr���^Z�͂�O��ը���V��y����܉/�6�j+n,�6��}%�X*���H�� ѵ�j3���,�RŮx�5G2?)�i��Wr��NC ���}��D˻?��������0gQ���I�� hw#�YVܸ����;ΨM�nQ{߿}����2p�ʘD�A��`o8���X'���z���5t�{�y����X�q)����M���4
���s(��b���	�ZCM�����E1Y4X�M�si�F��Dq����P���8$k)~�_4��$��w&�䀮5/���Px�@�3����N�3�`*���~�^(r���(վG�17�yr�%����\q>o:<�%���]���m�jo��r~�'&k��5'O]��CQh�&��~R��_�tƙ)��"��^<{0sHg�YTO(��� r_��@���o-B2Q6�u��H�r��+m:�1D*����%=Տn9�{�c���â�q0����E��� ����%>c��C�+���Rf07�zt��@�=������(d��u�:�h&�(�����0
F��z�_���>Q����QO�P+~d�Wgx�ȝ�=#�L���r�2k�6�n,X�eW��7�7��IJyv����nZ�R��@shN��v���?q��v�ϟh�A�i�N��<P�/���Mol��(J�A�C�/�t�D�X�G����;؞'�	�a�j MC�4�-�xNQ��kN]9�	Ȧc����H�_�7�n�Q�G��P#�зCOa�/�|��0�����j���m���*�u~$?���v���-Cٞ�'������]8�*7���܊���\�A�1��j�a�Q��E�c->5�/�e�8�j�c�����aW�Q�f.�.|�豏�Wm�gs��:T�������K����=�XW�C?�&��pXs�l�2��yŀ
���L�ݔ���'���AJ�$D��AՊm���яi��)+����"����q�9�a�q� �tݷ3e�W���H>��Q�@	!��3�bC��Q��9*5M�A��{/3_�T�[���*�3Qj��Ӂ��-�JQx�B\��u��
�'��O��̭v�M�/}�� �W7O�L�~�V�C�	�,6����.d�kM�뽗9���,���p�Wf!���[/��юPu�)"Pedn�t\(�~���b0  �s����נ�* ���?}��O��,��N�tE��f�`��}p����,�8eE�����޳i����/t�V�Aq	Z��n�j��Ac �����ET��֨�������+H��Y0�D���G��'�7�Ja8��<�G��^=��?�Q�i�*Oƪyˍ(!���!8��3_��oJ�$s#濕�.9I�449���fѩ��rb�#�[h9�ƻ���2I��3LW���o��J�����'"��A��??��\˘>lX�2������:�:���S���bznt��Ԣ� �'���R=��{�AoS�
ݗw)A`����=��A~,�&և���� �|�O�v��G6U��B��#o�c��{T ,�L��#�3$�6�ך-%wu:�t�Y�U�3�$�o6��y!8F��Ӽ90���ߓ@<����BL���tP�P]������Ni4�"v�ժW�2K �V�u{��Ԗ������x��q�ڀ����H��)4�C]ڵ6�_�W��ksk��Ѓ����c�*0=
�ae@'�\8 �7�ث�4�\w+�8æ	\w�}	��#��83�Pi$�l~�]���\ڊF<d��k����r�B��"퉵���Fs�Odm�(��������l�Fc�.)���5����\������O�ՙ�{�ฉoV�*"�_�0\*��B�t��7B���t��gƒ�,��4�M,Kc�˶ ��4ƕ�X�OI�w��ú(��V���<~�改�f.���`��Nsf�Y��9��>��hYr�u~�5x�/<����︜C#�^�Y����q��^��=�A\�*��3�=^˟Ϫ�) �,�V���n{>.W�{$TD��8+�QI�ˎU�ֹ��9��̀P#��mѓN�/R-ID#'�l�
�j���fj�� ������T����Wl��>g�����)�"q.+we���6O|��A���ټn]]Z%�%�~�b%���.�׆XM��B|>v4$).�Uzoq�˂��<�����aww��9�P�}s0�o�C����؁��ǟB;co=ۋ/ #�4N� �2�iɦ�:�A��E�Q�+eK.�%\�|�!'�1u�ۣB;�0�(���k{݆�;���6���.̯��uT\e�c��k@7�䅻S���-1ɯ�8�s�lF����������� �tQ�x\�c�h�������:�i��	�oG�L�G&��X�*��ɿ�$_wkt������꥽Y�r���4dC���n�ﱖB%���+h���t%ͥ";iC��Z/���B���p��O�N��oD��P8��Ϡ�D3~���YVX�M�Q`ԫ����C�g��eU�N��Y���ӝ�P�]^�6v�X��^��f���Nk�}
m/�ي{��@�a�F���	��,т�E,�4�3ZOn����!�;{����۴ϟ<���@�N��+���k,
�����O>��j�y~t�������9���qW�}��)�a#~(��Y�<��3��+��@ɕ7���BU���(X����=i��M����.?�_�z�3�n�N������X��ߪ���G��_�R�k�7h�%H�rT���'`4����Ϩ�᠁E���� �_� ���-N-F�L��N��6��4���ܤ4TD���	�Y����b�}v}�M��+�u,$�M��
��x�S�3o��2).�Kss����Qz.��V�/��^Sg&��Ic� ���7��9I�4��F^nϨr�p��6�T��q��NկQ�v��0[���'�"�j�O�J��DIg�Q5k��w��^���Cyr����Ѥ�{<��1�kk!b�E,Ѫ�{(~]'H��YEET�%��ͼ�d�K<\�\�3�XlR|��D�M>u�is��ܸ��,[c��h;>�e2S?�����qv ��+ul�؂��'���b��� E�o�U,�������:�Èx��EsX҆�z�^�!Ev�<��u_�����cbچ�*�!Xl�â�`N�I�Gz�y��		�7vz����6��1�:�>��ʺE��s��M5�i�D��;�^����k��a]?���d�R�H�hO�
%�S���6&��m����&�A/��K4�ɠ/gV����Ö���Ѥ@5��F�#�!�J�ty2�:�:�9���y��y�*����B�����|�K�b�Ѻ�v�A���OV������P��1��  7�A��IT*#��Fp�7�L
�h促S�g����%��u���i��!�k5��Q#��ah���V��-	��/��yĉ$ӝ��	��7���"y�����4V��_��e�Ln�#����t\�����>�����4�XV��V�`7k���r���'�G�4�*OՠY�E�6Dz*V�/E4u��:״�s�=���:Ne���{����a�d] ��6��?�_�]��~���x{&S2̴��e�վ� ���
��ݨ��v�O��
���Ƙ��/�W�h�'|ӕ���'{J=��K�PSL.=����V�3	�"n��^Uk m4^@kj�V�ʬ`�X_�j���:}��n��K��:��n ^"&��i�!G��#*�d-�(q��V��"ca�C7^�����6��ݒ"���ǘ"vh�5E)ɒ���5�8	g��B�q��,������!�І=�%��&�kz�����@�`=Z��Z���=��PW^�[$����a���X��½��>���wT3q�����|&(�u�����*�}P%R����Q�ߣ�j�b��+���QCTL/"���D�_Q>�������1��R�E��e�-�+�`S@%��+6�7{c����<�2�r��:us��N��ap��&��� ]�b��lV< ��� �>�G�X���ᓨ������3���QL�S4ci/��z����ۻ�m(ʧ�ܽfg�a���2�h&?PI�B�x�� �J	
�"5��4w	Z��>M���b�¤�>�fp���(N����j�C0���������%�c�zS}"F��4P&@���Nd��K4iKP&�j���J�%�������!�yo�r�p�%�-؏��Ȏ�M��@ $��!�E,"J��yH 0H>���@&8P9���V{�6ad$�f��δ�Q�88�&d[����?�8���E���ے&�Cin�,@�b����)6��V㴛@1X|t��f�9�=��e��?Q6D�$u�ZF�T������k3�!ؙr��W3�����:0��2�a��L�Kx����ѝ?�*��<��d4�|��^� �9���z�33A=��'&�c�T_��|eZu@��>��0�~XK������[��b��e����_N�
�T��Vv�;j�z�O�1�����������4(�yE��e�����' ��
F	�t��܂���ix�4�7��[f� }��w�<To�5��$p#��#E�8?�Y��`�\w;�ʹv�_2�I�v4�!�~��x�Jq�o)��s ��UB�Y�*��$8G�}��S+�����=?��-��P�f����+�_�n��|����}�S_�]z����g�쵳��k��tn#�o5a�S,q��:^���v��
�0;����ipo*�T8�N�l1����6U�G;�B�y�oj��nY��	&����*�l(��=K���:��1>L����A��[�Ԭ�d�0~���E�#B�a��F�`��a�x��.N|�[��Μ5T�g��-�_�a������������Z�PBa����.?�k �Y�U^��=*����3y�FZ0UN+y����"n�g'��=��5OҤ����ᵨ�{��[������2?�����%Α���ƙ������^���B$�o�!<h�W��eʈ7�����0����{pg%W/_K!y-An�j���D�)�4��^���Z�������=�e��F�h7� ǣB�JܛT�_�k��H�	?>@�Kd����U����cR!������G&�����i�����H1>�j��{I� C(�C� MD	�GK���0>�ʬ�ɦ�k�)�$ X-���>|�~�ǅN��L�܄�<`s�'�NQ%,[�Ɗ����[TW���oDa@6\y����6��Q�`�֤�ET=�ұ����a8��t�0Cg&��Oa!�2݇�Z�P��H!��k�Lk1|zA&N��U�H��Y�	6*�M��N��vD����L��u��_�^)F���B����8l@�������_HWE9�fU)���l#R�SH�34x���c�A�ir�\/��,���B���R��k�G/�t�KX4b�]�Qd� �K�]���0]&M�H1�xA9q��Y�.W
���n皽�X��E�&�B��|���7�zm�2�����@�k�/�R ���[�S�t4!?��2�|&���|]?
�:!�1t��hl)@�a���<5ElwdT�n����\L��T�2K��Mz���@��J!4m�d�;�}��)�^��8D�����cg����_G��Xb�����\�`���x]7�殓HdІ�fM1����B�z�>H����7�_<
�b��U,�/f���?���t�{F4���n d��{A��М(�}}�y���P�d����h�KMU����4AH3o�´]���������|K���~��2�r�y��mrM:�
j�����,#8R�ؙ�zQ���BӍ��ml�wq��m|���h�״oJ��f��*|hg����2>������-���ɑ᨝�TD0�9"�PZ��%`~�ÇXW�%'G���D�0�ܦ��*�~�0��l���X��XW͕��$�WE�\����We�8��/���4�ٓ�0�6p����v�(��;�yA$'}h�P"+ ��:�����u�����d�3�*i
B.*Y�Q!r�6IVo�[#�x���8Om�8�Ƶ�g\Օ��[��C.έ�q�DF�؄�&��1�J��T��P�3�@��wÃ�UC�S�^[;|��1��5����a@�'��vf�r��Qa�H��|��
����$�E�5���Q�q5��=�e���z��@����G���)�ns0z�Y�e�,�8tA�_�7�%\s���]mFuR���­1j+]{������d�q�<i�#Y�����ml?E���u[�������X��J���T"h|D��{�jх{��G���ֈO�Z��$��ɾ�C_΢@+d���>� ���҂�uFX�A
�;#���Z�?D�r޵����#�X���1}��K0D0��N��m%RU�*�I�%��S{�������1s�g0�i�����*<4;����?�#�?�۵�+��/�LOj�����S�.T��)�/�g3B4�d�%�W(��l��������Ze�N��lKO�yv�����)]+w_G?uC���s���uz��)���8z�X�%9�v����Bˊ�	��I�VE`���`g�2�ؐ�ҷQ�C��Zy�
�r�EK�M͚�x�e
Ȇ��e���A��+�?c���l$r8�A�#<� �S&�.�u6�M����>;K_�s�JْX�fYF�n�`����,����O�#�Zȥ�8�(�Tҋpo޵�$��=�g1���u'~Zo,���U
���c֝�|z�s�A�t��������	���P�A�i9wy7�Z��o���ؼ'�s�P���t�x= ��l�Yt ��os,�޴J>�9و<�0�h.��C�k�T����-��f
�M*�&�ٵ�?�W�PA�
��wձ����������'��,o���a��ɿ:�s�Ljk;���z>�mb�K��)�h&-qWN�����HkvD�ٰ=D��TAk�c"�#�'��m���4aEoG|	>�n�K�;D*4�ʢ��cCZ���~Y4?W��U��B(����)����]��9"M�|���qVH`�I���:'����⸎* T�E�^|0�Yo��m�J����΋
�:��p��w�V:����\�ߖ$�ʴ�t�d�ϼx� S���B�CD@�Ԩuݎ�5�B�/ρ>`W1��94]����R?,%Z��z���(VL�m ��L���9�,cw���
d,5�U�D1�ţ�3�(���E�e���� _��nM&!\.\4'�>
ؒa�P�G�lOM�n���] '��K�m�,RAV����^��H���g���N��ܓS�klN�m� �)EP�ׯ7{`�nKy���^@�r�_´F\�(@����Cvrk#>c��i}�X���]��Za�h�?���0GӢ-�%IJ%������|�Q�P !�DY��P�@��s�%�զpl�綎�OΖ=�F	��B�������U-/�]b#���ާ
zmU�з���Ǐ.�K}�ݧ����]�P��Ru��cK�
*2���x�a���������T�7���do��l6!3���*�o\��
��qMdm&�1��K�������iq�|����b�ce��'���f�,q�k9�>�� ����� ��H��7�H-╟+���9�k�uI��+���k,���Q�ظ�zs?O|��7��/_�cS��=�E�j�Ѐ]��˥��~i��<Oxs�Ѫ�1�3� -��9�I�q�{�-�)��nL�����X4�Nv=���}[�WckO.��'���X����̔G�ì�4o�*u'��j:j��Tj�!�f[*��# �������߉6{ý�d�Ht�I�Y� ����fN�r�gi�go� J�@�\��ɐ��6�3��Ò�$��*�!0��O�I�'ߣ�[�f�&�B�]���I��'6q� zaw�t��2]�����`��|�� \�E���4V�a�+��j�Ur�.X�j8K|2�E���l�=n�Z}&]K.�[5_.�����чp��5�lٓj&��@�Ahb���w���\y]j����&%Wk����Fsv��:�~:�[b���{��Η���<w�-�	.F�VRQ���1mWd�3��@���X�O^����/�97;n��*;���4�R5��v���!�B��j�?���_����7�e??��=���7��}ϵuˀC��!B�W�װ-7�H5Q}L\y��Ӂ��]���m�z�6<��0��ҷ��� l�ap?(Lt;���E��ؿL��J!�����;��;l �
�S���v��^g;�dDz*����fh����U�]\��~�hG\#|7Pos��4B���Q����|��v�=r�&!L`��5D=���u�n=�Ltu��dP�2B�0��J�-���L)WK (�7���P�Q����'��.b�ˑ��	�R�|��K�$1��X�=O��(ny=�sm�UNw�D����*�1d�e��%qT�t�
R��mf�������,����\���2#�RMp�b��%�C�����	9�� �����5�lk%<V��#������fb�f*��Έ�l�Ap"�hh���y?IS6�� �{�3{��g�<�hgB�{��#�YN(��|ר[�gR�K�˲>�hy[H�z?������J����月�i�Siu<�c۱�EQ���|�ͺ9�a-
06�~�����B����e��	��u�(Y���6�|���إ��e]T���$;����9�(=��X����]�6?n��?+WUl�@@�=|����Y�ia��?J(,�$�C����y�22[�S������Q�C7���<�5z�b�.�,+K��V���0	�22R�Ecoե���K`�|g�3s>��-p%Ņ���柪���+��:�{�TWV�|Ɨ��W�A5�y�5�b#�D��{�PY z
��A:��>2����u�Y1IO*��R�w����B:��,���d�q���>	�F�����:��鏉&�����)X����?������=��Q�>�}栃��A����+h=)�X'8@���^6���z�_|A0���`��ס�)��4�gB� �Z�9x!t���=�������D�|�q�,=3(��@+>2ۚ�?�~M,N�K����]�tĥ�sy��*_�*���T���f�E' dW��w�M<��QU��h-��?���ob�.���Aۨ"���EbҠ\�&����tF,8=�9O6��?I+.md_���� ����!�����M,�6��g��.�UK6&�9�_I[��bY@vo��Z΀��X���`�vc,�&ݧ�\"HP����!�{u{��#��t$/��!�p��u-׷_6��hM�P�24{/Z�5�L�����?�#��7�+N�!�sk�6�i8np�X�M����d�K������5�6�����3�ϒ��ý#��.hV��|�`]�=�+]ｇ$�y�fuU?4|�Px�NLo[*�:cms�S�Qp)4�t��h�� f�@���V�"}��Y��L<�H��g��x���`	�jsݼ?���5[�Z|U�+0�����C�6��!�+?Տ^�z?�����niaH�^��)vz��)أ�6c��U�{./�⶗x�{
�h��2K�ޘ�S7�I �iD�2;�Yc�1yׄ�BL7ذzz�'�J�Y�q��;\\C�7H�i��8K?��{�R�ƲhԎ�������yX�\.3�C��6�͚I�N��SY���F~�E�>?)�Vt8��4�Y��7�����W' }�*/
!�QP����spC�X�\q��;1������ẩ4�'i#��eᝨ�|��rGn���3wKWb��*b}��f��M��s�4ư�j0�U�j ��%_>~��A '�!H�B0����+r��l������;��Yu�;�H�CVt�Z1
�����ϟ�G��?t[ae��6GCZY�������EB��BN�_/12
�w��#p~+x��{]�`?+�g��В,d���8�mt(�TS�3C�V#� ��֧rF�Kh��#Z�C����
����吶7cHbU�R��EX��F5��kҹ�߸��)�`�B�i ��uo���̍i�O36�pH��RQ:k��a��u�����UkT�[l<eK��Y���C�6:�?wV� �0B�^$�������zM�nb���67G�t:��O����������o^P�ZV�A���� ߑ����OPŅ���R\'{:�ſ�Fݥ���#�����qv��CIڵ���@�_��@�ǝ���.Q��V�|#��y��ϟ���#���>9s���Wd�1W:�$���j���
 I(�mW�#C-Z�}n��u��iڌ�N�3��?���: Z>X��9�'��[�l��L/b������A
�%`�=�HO��o`(�MR`�!����NI����y �/,N�s�����Q�x�^��[~O����и�@Ӛ��5���S�tS)�'�q�]�f�T��j�>~w��昔���a"���rW��:��7���3��W�{E�Q�:uTJ�ka��'7E����XOk�;�N���B��X�V�"�c�Q� �lHT�����#�+���blOWL�Ew��Rn���g^��W+״�r�)!���A/�/�#��)����<�j%�����X\Ǚ"hևx�0%J	����	��t*�CUR!�hÑ���Nh��Ս�A���҈j%�٥�|���o$S��\Z鲇ڢ/z]�zXd`�h��ĭZR0�N��E/����G���vqLU����{_�F<��-���%�f2��ugz ��3: ���n&��5I�545����H��ye�hÒp�ܙ��N��\����rr�l��t�Z�����ŵ�0���|xL�z���x�`Ep�3>U�ĉ}j��,�W^�18j��Q\!`��I�$a�h1o)9G���1��:��Dv=�[���z�MO�J�۠�
��ׅW\[����
h�����Xӡ*�4{�b����d��ͲИ���\WT��\mʕ,9��P�0�AP�5Z}��ר��^�����+�;ۑ�ꅐ���fp��f�T�,K�����c�{QF3\G�9K���cE���$v��à�]��TB�m@Ɋqw�D~/�sR6�y����r~ۃ�7��ȶ�3���/'PTu�I[��֛�m+�+`4�W�B^�5K�0��d�Ze��!v���^f�XN%�+6���Xo�7ڲ���4.T���.c�{��cI瀛�ԟF�b��=ӵq���D�?#�R��/g����@/X�	5QB10��Bc�)��Z���E��9��NA$��N�+R����"�w��,1֚m��'�b&.NyH9��y�( !]=��p���L�rw�(ټPc�V�UӉ-C�+5�B��갛4q��"�,˕�`_W"�
1脻X�җ�X_�kJk�TrVOs �/��wl�EU&��&L����E)���.b-/�'��9���S���#z�j���I$6OR}��Q�$t��5�3H�<�����%�oC�ї���co�g�C�� c� ��%���y8#R�������R>Qݧ�()��w]�����+��2�.ld+8�eĎ�&r�4cau�v����)Td�l�{�����>��nA�i�љ`G�W8��(�ū���J�����f�3�@�8����:��805{3���1c�����kq�a�\j�Q��j,��aWx^�@>3(nJ-��ӵ���XH��gͮ �:��t�\)���clT������*�(E��ov���ch��e��`@�]"�ռ��|��*/2/��`<:94��h_�&�r:p����e+�H��<-����sm��t�y�gCXHR���/KQU�
���v��@��1���zӀ^m@4��L�J2*q]��7��|,�u2Ƥ�d�u�\���Awݡ�#{����,��մ '���VjwɁ��éJ�H��0�PX�e� t������|�#cm9���e�A�u��p"���p�(��a��"�2��Ⱥ]�^n����^��p���/|-�"��D�F�_�$��،~	�N륱�����\Wp~����}�֛��Iǘd`�����v�<C�]KU�(��)ǙD��R�Ս�����<駑��u@a4��M�XO 7C�h
RD�ޅ��?WW��b��L�M"/��a Ҧ͓��[J�F�k5 9p0���#�ϋi�EC�;sԘ^�?��D!Y�0	�9��;�nR ܠ��A[r>yM\(+fL�3T�c������a㾝RR�C�X���Q��N:��W:y�zq��Ŋ�Ub߷���F��~����h�Ǧ���iu��1�g-��*�d`�6ZYqv8@�Bg����g�G n!ƏT��b�]���8>ii&D�$*�&��E�鄦Q8<�Vu|}8��2cc�z}fp��cMM�{~N����;�����p��)�f֫.ϴ� E��L|�T����m�?B&z�õv6"3�����ۏ.Q��	;��׿R��4
軍�P��@,��0I�F���|Ҕ�rxį���*��끉{�OΟ�-�')�p� �R����UJ�<5�O4��z+he���˽4�q��l��&��%�{7`-�@h��wC ��� �7A��b�0ER���Z�?	fM�{��}�f<"�c,m�Ȯ}qތp`(_��e�zH���m �O�TV�Nю��W�x���v8�c>1�P`���wo��?^���O�=Z<�t�t�6���UM%�Ȧ!|� ���J)�]p�tj�K�&�W }�5=p=�I�qï�%9/_�ﱃ_�%$tJzǎ��ĵ����5�ۻk���߲�v��1ۇ`
�Rٗ(���Z�>"_�>}��X�+��X�vߕEtÉTe0�y,�m�y!�*�Mr=�P t���l��n��o��F�;J0-�*N�2�����2&��c����@�R��³�l�8���h�vIhɞϔ�z��u����~�
E�x�?�X�օ�$���K)�n ���p0Ħ$&s�4� ��O�G�j�� (1C���?NDL�#CyQ���)�p_]��e����f'H���zy�xh���(X��p� �4�ZՈ>�ZLH�09\�F��������9�%�h�W��A�1�`�3���^nD]��{�G��Cu�fr�58���]�(#x�/b8λ���ȴ�E�\r��
�I#ʆ91?)5,��-yejg�Z��N�9�5���ۏQ�����:�r�g����~U��ML�F��H[0�L+�����+2UWri�IG�|�@�E��
f�Y_����g��U���c��u^�����hn��3T5�o��x�=3v&�! �>p�p����Pk�v�+�[eb~��F�����R1��S�"���*jc��7[@.�{��
�i�s���Ǔ5�f͒0�_65��06>�̴�Vt��h�c��������5I�ô��ůd�=�t�35���7w���nݹ���w����Tп�ȣ�<���5�n%�W��m��D���ИEF�D��6H�,d��'���c��W=}�Dcq:�9�m�p�������#�2�'���'@�$6��������H���PHB�C�V����92�N4Z��;� ���H ����jU�w��^���8�>eS%�X&��"_��E���Hq�d��n'�����c=�g5X������~!���nQL�Ҧ3�6�f�y���#��b��L��
*HDm=:����lno^�����_�<����#���Y�UT�}A5-F%W��ZY�s���9Β
����G�*C��fw2����e���gE�2c�	+gs��P�VvK2m³�T9`A*���Iր/M���I�����g����M�K��"��nwxA�)�㐁�[�S|d��eEg���t��6|�W{�
��~���P�ݠ�l��$;�݅�
�������lXo���aQ�[vÑZ`�S\�2<|Н��ҋ��+LF�V�_�Eȃm,�tu��`�f����Ɵ���ҩ�'6��s\t���D5�мV|��EJK#�f��Lw�$��"�/;�S���&�d����hĹ<�W7��vb[D�I�6Đ�XE��+ڦ�lP؅��ݨ~�P��	@��:C��=��ԍ^9��T�&!'��Ϣ������e�AK�VL��L'՝xK>O-���
M2	�t�qvj�Z7JӨ�L�J��=*}�ћ����2�.�������~�ڤA�}{���,� -2S���12[���~\�A�����(>�ܬ6]M��Z�k�o�9��|�������E����1����$�GY� "U���ծ��X\���+օX��+�J�'��x2�������>��9�Ӂ �F�D�^��5JA0�@�i�-E�J�B�p�%җ9(�P����m�������rM�IT����d*�����\�Zk���.������φ+�9�Έ��<�y���]+��g��-�ZQZ�;���=�C�����t�&� (�[��`����oP�q�ېü���x��P�K��%��Zΰ�X��9���p�3�����ߐ�
�I��͠�\���������X�ȉ%�0�x_6n�nG�Xm5��#�1��f�2�y;kV��\�kk04�^'k����G.�pg޲�L��N_%g�:�֒���zq�3B��d$�ϖ�����[��4J	Kk�HU��K�dy�mcq������I];�f$~#r�Ș3Œ���Il��|����9�nEM^R�#�oܕz��@��]�������UO�l�������`��5m���n�%��1�͢���Y��%��&z����wXEо���prĎ���	ϊym~�:|a�qto���N��Xev�RdOR����7W������~�km==���~�P*��H�e��nYg	u�=����Qک�q���v\�����n�z�BP�t ~���n���UY�?�O��{F��8+.Df�f,�I{7V-Z݀�y������W�Ԛ��
����=8g&��*{cR-�o�"7�Fu.-Ctد>��]-��Sd2���$�N�^hX�V�3.Rt#�B�6њ�@$R^^_u
We(����7{M�mO(o�Ι���`���W=jw���n4��s�U5'	�๻-���=�C�~�A	Y�����B/7��O��H��P}���u�Ga5��C��3�{63��|q,�W�I-A	!�.!�4������z����{^A�c|�qZm��K�Af$��-f�g)"� �r���D2 ��$��Q��U����9�&�fo�k�4��'��s���H��l�������f��9os�4:0?���e�g�U)}{�`3� �����
}����I�Z�� �|[!�$�_F�A^�E��D=��lK�Y�.S�۳��?@�}��n�9۩f�� e��"M��`ݥD�|Y��������[K���u����Ⱥh���i���x(I����&I��;�dj6�Z�TM�d�sh�qT�i_�0{�Lʧ5+g(����N�����`
f`K�! ���Tk��f��E�_P����@����vP@�Nqw��h;�)~2�J�$��!������ �w{c���i	�Ú��\�ܭ=��/�ډ�g7l�Jd�;�Z �<}��y"d��t�M<�q�i�2\1��Л�w���� Ή\�'��u
�EHִh�V*Mϓ�O���`��Á;�B�b��U�� a��:	�"Vobf�@B��S���M��z��ZgG�������y�d�s�
�(�g�km�@�R�+�\�4~c�����b��S�_���/�v�7ڏsb�'Q�U�����]R秷��Y�Kj	$������V���x�a�q˽g�Rܤm}{��GO��`��57��0pr���Ś\Y��slzgG���lRY��U1��?R8���h��*��T~V�׹�G�j%���o��l!Hn��]A�4�Uͳ}����bfa������;q�R�@m��򛧥N�!cQ�|" ��{�V�r�\��H��Z�7~ǥ$����X�8���wꮔ{T�$��SV���������5�e�u\J9�{��|��M
KOw�@��G�v��F\���d�n��_������}�i��=.}]�e��Fؘ�,�wlR��U��hUG`���t��!���`����~���NP��+� V���{C��l��6,��2�FC+�@�~�ؓ��	yn�l�7�zʄ/��n�"
�<ǉ����4���|� V}z���F�\��V�P���l�!>��s��&�P�򜚁�%��5����*�R3�;7�`ZoIU.�C)�Ss�?)*@�=j?5���� �剐[q.X�v�-9��3rF'8���_b7�ۚ�dIp���Ԫ� 3Z��0r���:V�i��n1��r2�|l�A�"#4<5��OVF�w�שMz�j��y6�7��ڊEY����21�(���#��Y�C�恶/���=y:慖?�/�g�p��깥U�ފ�g�HY;��X�{�`:H��u�5R���4���&,MM��J�13��N6�.xs6�6��-�YH��]pc&��/[�j�e俺��w�u�d���S��)Ab�@vW3&��R�۾�V6Z2��JI��"�;�|S���S�/ss���m.�wxml��_e��n�1��%�����Y���)H�ٶ�YL�P��9����I딁	���d�q��O/<�S�HK�Yi%�@'�S/�S~u�x[�B����!f�4�s���]i|e���1�xZF�2,�C��'��ҝg��̭��
X�D��S�P%^�$j�ǣ_p�z�ԙ�����V��_�;u᧒T�R��em��m���5%�9�%�7e���>~�2��;�/�H�uj�/��~���/,`�!"ob>|�3ꔋ�O��!R#��ٹsJڤ{R��-��H������(|��/��t+9�#�D����
�z�.��u� 8�
L���\.��Bo�~̄��ݎ{����2N,-��[H:y�>��S{d��ۛ����ܑ�Si $q�_"���N���A�3��7��ɹ�o���wc����d��Wm���L��?�]�-u���&��*{K�6�a�#G�P���WZ���a+Y�FN0|D/��Ȋ�S��k�U@ �)��[��-p�,�C��ʄz�Bc̅IA��O-s���.��I���������;��A�%�����-�#g?"���17Q\1��9�r��
@f�o��~:9b>�����|���x��l�Z��5���ٓ����\��Fa��������q�YG�:�(�Uĕ7�C�P��ug�9]���K֗Ei��5��4r����u5�Eb�ѣ�l^F��Ҥ�0ev\�xlVG����7�����-v-�х��͂i&�?rc2B� ')=pg�S���$H���`��\cQ&P��� ��ͮ�i��v����S$��*לk����'#=��2�wU5��o�q�3#��w��{h��fwJ��t�҈l�4a-Xx�����Ү'2�c�G;Z�+P�5DmC�������n�7q*(���t�.�� �T���E7M�蛁_x�M����9�7^l�}�"��;�q���7�nF��׾b%��%����!��3{Sb�팃��-|W��.�R���;�NNǒ3'wǞeYYy6���Q�.3�X����5���=~��H@n�p�7쪙7��xo_��W�ۓ��d��baK-E�7������⤕��	[XZ�0��n[<A`~Hm@[ �ꭶ��0$>��)!�	<�2�� �[ޘ��̥���B�x�f��q�C��=}��LP*�.}4�{A�y�?q�y��-k��������D���w��Ds5�� @�.jJ�H�MM�������?�l^����{zET.��/�Kjq�8#�3hBEq"�`�P\lYu��KG딃�g���������<��U����3qS��l54{�}pvh�9}G��S&��3� �Gx�o�ӷTXQ�6�$��/E��&|�*�����q�C�=%���5���"�%��~V����Y�ئ� !��k�8?��75�ִ�o�z�(���2�an�m����t�]���-?as`����g�h�xn	�\�="��C���4ep�j]N� !�T˴���i������,�~�u��e�{	ؗ�-l�oК�b8��)�ف��p�J��M�%�.ٗ�X��P���n�N���gq�9)a��7������e��x�iX�����Y�����y�q�D�����UuX�?C�Hń�A�,��*]'�v��^�S���/
�3
.�Y��zV��`�%�|<dW��XZzsus(|�`.jY�Rf&��2��aR�#��T�"(ݵnJ}���h:����2��!��A�>Z5����N	��0U�1
��h���,`�Bjx��ԆӈU*��7;���,�]ؼƆ���9�� �^�+~PA��%G��Ś1t�7�+e7p�L��b�	�V�-
5��U��|�M����Y�Z��=��hYS#�X���	��U��,̯3�bd��:��B��k��$Y��AVtx@(������Kj�eɤ!eo~��Fa4-ŎK}��PR�;��|��M���O�F����-Q����%
e@���?y�7X�k���a��H�7���-����^��Ί;wln�Dm�����^��*�O�m�o��������UG?K7�8��C It��s#`k��.b��:�Shoq�̮�<	����EX�3:�	_rD���f�f�$[��9��WWSN�XqEMt:5�}4�'�k`ސ�����t�R�����s�q.G��7\��K��af�Ę^m���ɾ�R�ːB|�"��
�/F�3)�*���9
D�|~;絪����1�j	3�΍N4��m^gժ�v6���յ�'r�[q�5e����V�2?�&��d�!�G{䤛�4��'�zr�.�R��B&c�H��`9��%�$�0���Q@����t��i��rT�@����ް����S�-Q3�?�Jv�
�@~t��O)��2o3��^?a�Z[]U�v�@7>C�9xv$Y�X˵&�A�Ϝ���wI�ϡ�]�'�S�պ�l:���V�RHB���M��D��J��k��
P�I�ǵq�}�����	`| ��Zo�ͦJ;q�t� /[:�*Nm5�*��L�:�x�%n��"}>l�c���k�"`� ��>Յ��#�\����WN-�4Y�|/M{�OI��u�Q��K\���]�hT/w��!�m�]�yF_dL����7t��س�����s�Ssԩ����q�)>�EЄS_�Ab����Hk7_�#����P��S��(�a��Ovx� �/�4���c��6�)�cƷ���}໗�V��*�H`uħ1�4���	�)Բ�]%�F�?s�S��U��{�B��y��U������{�JW�Aw��o�jg�ۤ��F��H�[M��_s
q3�־�y�ԍ�K��LS1J��7�M�q2��F|y���Zb��O�D;��د����E'��4]`�l0뉌<�.�g[�H���\�/*���\y:3�Q#�׵��C@\z��s!�)%�"K��{AŃ>��K|��<O|1<��
�P"y��1�\�$,��W��C�7�؇�ZNb��U:S���`�]�M�J���1�@�fz ��^X���$�C��D.Ky��o�hlr=݂�B*�BWv}�e�n�RC��,��%�F8'u^�x���[�йM�qV�FG��ϻ�țSk*D�j�+�?��k@k���Y�Bw�f /�i+�'x�M-��t��k㢚���r��S+7�ײdъ�j�����)c�h�\��EP��M4�bC
l��(n	��;�������\�{ƙ-f�$�lǗq,�8�[����T4������N#�	����;�Jj[Z���_��'g�v:��4<�����b�3j��m''�=������Y�(`#
f�R�b��Ƈ��Yn�����v�&=��c�_:k�,֔�u&�~���'��]�o4�Z���u��8'�	=!�V��(���M��	�
q�>ܒ߫�����̈�i�e61k��)[�+�v�vb���$�?x�t�0kq d�$vդ���s0��Dm8�$س������!�ƅ��ö�
�B���Rd�}�X<r�oȥk;f���*�FQ�8a�d1������&>�o��]*�Ё
h.F��0ۥ��{""�_�%�G`^�:n���`@ᓷ�S&x�ٟOH�y����0��|;ob����Ma����ڰ��9�e�]u=���
��Y7�l�5��E��H��R���b��t�d~������;��me'�lh�雜�Pqyt\q�/�c(��}C��Z�k(�(�$mn����o�4�2���U_6H��L׸`����]��hF\b���eٴ��X����&ԅ P<��?2`	��kh)�1B�yCn���(~��e�s��?4�U�Vکㇰh�������9(���]�y��Do��� ��	U��U�?��ς���t��
Nn�I��UaJ�����3M�xW�忴@�ב[��ҹQ �x<EQ���1�=,�mo�s�.�����^��]��d!R$椌�#�K�I}Ļw`N̳I~���C�oS�^H�:<��v����q*Y��~]2d��Wq��e)�>�􅏼�����>k�ᙊy�6�[g&�j��)H?�د����{��G�f�Bn�;D,��d/WR��N��L��)�����µ!6�lV��cV�*��H��6wKp�"��%Q�4	2$:!q h������Z>��.�x|e����f&\�H6�����;�T��K��T���=I��"_IO��J��X�*).i��q!;�1�<MD:��޸�FGpv��e?ݔb�0���[��������O6�������Ai��KE��\'r��˨�w%�29���J�6�`�*���B���V݁�p���_
ʗ��k5��	PS������Rb�_ŭ%��ܟ窳�-S:��"m��JU�ϯ;��c��C�r빞	m��ЈŚ�IS����c/�3���-�i���"�A�	l� {��e�Z�g�q84���a4+3�q��4�\y=�of�f<ւG�%���P�[�ý�g��翇!�>�{/��2��! �lD̀�9���o����~?m�=��� ��.��U�j�h�az({��	��-���7�����H���#J{!�y;8��t ������{9�d��9Ik#"pq����k�Tv�Y��,�NÈ�{ˣ�pG�<y�1�I�	���2���b�
�@�{_l��Os��e}2>��d�K���Y!cVn��@t+���v�@��S��E�o�}��*��-��P:s��?x�tĪ!�Sk]Nw���7Kϒ5pj��N�k�{}�=�Y�M:�jo�v���P��@z0+dN"�WZ[�����"AcLh>n���r\�[���b�<���-Ø
`�
_vz���@�>B�ZЦI�B�	d��c��?�>~JO��dp�m�����Y��J��Z괿P�4:|T�D�e��1��GW�$���:�*�҈���rtk>EDˊk�o�,�Y��%61wT��'�0�a���/���\��q���G�a��GSh�2��-�7���D���ϳ7�U�?�~sіM�e��t�':�s��"A�!T������{�N�!�4�|
e���[��fg`a�eoR��iZ�4�p�^�<�I#ٱ#��&�
�@S`�N�T�D�r�!�#*A�n�S�Mt�yL/�u�qsQ��/�a1�q8�DY���OZ�i^������Y��4T��g0�/%��y+���;���w���� �k�=��Z��O�N�)"�Q~�8�g�QE��t���G�I��x��Бip���铪Y/pi�\>���P��������o�w�<��9e� igv�:V���ݟ��5��|Ѯy��gj�Dz��q�����y�M4�'Y%�0��)ik���5p��(*2{b�&�-Eq��cg�U�F�K(U��4΢`��I_���>�%���ٮ_���;�����j�; ~��=dn���Ζ47�x��3�ZS=���^6�������jE+���Sb��>�\�-&.�KmS�	(ņ���f���ȜQ�����"�u��EaY�wC�2�hҳ�*	�-�\�p/,�wv$G�v��Ϲ�0��K�x��L_v��ϻ���	��n=c�\�s�t�7�K�Ah"�~�8���\-@���`I�~q}g��dcQ�_�Jc��V�E6����	'��}���dxqC�g�:�����R��7P��܏h����<��ڟ�r�����$S�F��1�vh��%�������w'Պ,#`3��3�;����C(�H�,N��,����Y���Z�2#��i��qp�s�~Gq�8�G�s'�P<�6ο�2
�^Y��{#�!�l?K� *��r *���-�}�j$x7�ɴ Q�r�2i�j/a�a��h�����׬T}���@.u�ǂ�d��b�*&���ӏ=W8����4�N�o������zd�n�GĤ�C0CV��!����/��U���/�������%Y> ���L�����c0�I՞�U5����9U
aҿp��}_�v� e��_2�4�	�]���jK|^���g�NV��a޸��`![�5�j0�0��Wd�S��<�͊'BG�N�t�"h�Z�g�� ��VO�ڲh��n$�F���k4Hj���\$f��fc@7)�1��9�ԋK�\c��9��ؓ5L��K�8_/�[2���'mhK�a0��"�r	M�=��cH����� �OH��E�����*.0�w�o=�UM�+��J��_a�#�
�to�Q��|52�H���{�Z�s�k�Ƽ~������%�ܲ$�]�A����+j)l0�M���H$��~5`���iPГ�3hO9~����&��*��DЫ FfsB�r#w��[`�$gH+lvC�J�������U�c.qB�� ;9l�e���o�x�|~���Wѫ�O@��F����O�F0��1�Ug��U�J���8%w���T�1���f�K�]t���3�!��� ��q��ѩr��/���~���L���r�wP���;ODvĆR���K��)��ogڟ�ؾ�$���B����P�\3=S�B.�����r7�%�����F�#�=���n��2��{���B7�"@s�j���T� LfzM�I�gi�TU]V�����p���H1�&���t�a�w�ĄFW�j�ڔ�4V8��;jc�<gCT�f*����lAˏ���o�[�f2چw�RY�Y�r�b�xg������;��6�$θ�%_Sf� a�5yp��8�8��9b�	A.B;a�n?O�N���M�Y�Tl���8t�屫�Oq��&�S�"�d|��X�ʂ�{6F��'��6����@�Oxt�ϡ�7�g�Fظis#���FK����"cY��%ޑ�~��)�����dx�����b�@�\�G��	�#�$���b��X���Z� ^ v��l�o{U�^����zM�w��+9�氚��;��/�ḿ��6���@u�+P&��]R�?�<%�M��,�Y�v�SX���������k���l����ur��M�%���k�a�S8W=dL�<=�>dg��#^�:�����uq���Be�����-���;�B���	������r&&���~�t�1w�ͪ 8�C[#�@�6���SS�<��.$�܎��;v[o�.���U��V�i%6�g��ݮ
T��.�R� ����hd�?ܿ�oԫ��i�H�e��s�R	�A?��6�hT��u��'�yI@�r�:��8H���?����7Z��GUH��<q�QD4	��}�i^B������E7)��1KSGMٕ��ɔ!I�������C���Œ:	j~_��ł�ס"�9��v`��,�MݽQu߉B��A��O\�>;ٍ9�nW�*0�9�}(&��~\XS.�}>e���k:l���:O�謨#�7�~Q�C<M�s��������e���}��P�a���z�cZ֦0���Uf{��W������1��[T�)�Oni�4��<�S�-�]s`Nf@/����v-Ȭ��V��^[�����+Nst��H��-����Xx�g��Uޅ��ss�J���ZW�4V'��Y�g̧?��W��ݢK�)�O��s�/�;�~��A���Z+Tۺ���'LDNuBK&!�z+��1^��9}��rfqi��t�k�D���,
�N~�Yv^5}��C"��� �Y�ρ3z�Gn#T��\��%-���������!����!	�y��]��_�.N7��*�ՓuN�;�>�"���D��m��F��_A"觠�6�cF�ea��N,�!���"��P�W;^�4�̟��{4�$�Բ ���b�Q�D��ضá�^�ّ�_� ����� #���W��.��9~=�X��I,F�;^`'�1ɗ j�5X�Xo~?]E�)� ]��1~�q����W)�<����*�h���b�n����>����x���-\�~]gdN�T�G{�{�s���uER��H��\J打�V��(V�'�J?�g`��%���e��P� O�!������N@�Њ� d����$ܰ���Č[���5_�i3ܖY	3�"p��ۙ��܉��|��qÅ��9˼�__x��%�z/����� ,�9RP�7�-;�v�}���h�>m�A](	B� m�fg.i�}K=�]��ۊ��xfP�z#��4����S��>�L;��M�:F�LaV7�6�1�JM�B��uj;AFO"+��[�����<,���F&�b���M���6�&'��`�W�+���/@�/�M@�³���^[Or�?,*���'.r����f� U�+�y3}�Ȩ��r�w�q��$
2z���4��e��$��k����[`Ψϛ��mΛ.AH%M�Ĕ�/��݋���$���P�+���~
���p�	[�M������`�y>5������փ�W�+n�g=oMC�"C�	�YS�ϊ1���B"b������k�R۾�ʕQ����p�f[EJ��O?����/��9�/�ؠwr��<�Nj��շq�őA0��g��]5�@r_���l��a.�@*����2KN���Z�����$ ��H�z�oH_p�dê+z�Z;a�w�Ou��7���	<�2zo.M-�~�ǝLH�@����޺)�u��0:�/$qOvГݺ��j7�gn����=�2��]^'z͓N`['���'_�AFVf�j3[��z\J.�@Z�a���x�zv�,ǯS���%�b3��ql�<��B�2h�e���N"e!��^��F�S��ت'.�&���*�l�8��`@�'�G����*1.atF+�^)�Q*�&!�K�X�p>��I_�pv	�?�U���{���Z�p|Y�Z?BS���'���U� HQ������#?��M���*�)�u�1z��I��.Za���b����B�ר6x�9���l���O"�ܚ�l򒍜w�:�$����Mp���E 燭��ʘ-ȏ���#���=f(V��O���s\�QE�?=��PxP2R�%]R�s�7�d	/y��5W<6���ေA460� �U�C����L��h?�k�5��$��>D��� M�p�ȇ5�a<N��X3n}t-��	mh}�V)�|�+2�Bn�;�D7~Y�E��/Na���}�)u��5t[��p���8:̐���J	u৭ł�U6�\|M�z���)��eL� ����1?X�|��0;o���dshf^�=�I��p%֢ճ�yӻl%:�!o�@oZ�|���.��=�y���*�Z��|֟��}3xmnR'��p%�X��]z]X�e��m9l������)��G��+��3P��%,UC8�#ݬ��'�����C�P�a��	�.�q�1oL�����#E�ِ�}&��aYn����N�T+G�E���d����	�1�T3�(��s���ŵ�z �<��G����s]�R����B	���&Wg�D-qS;�	�]=�k_��M�)���"�@�հ�'QX��6U�-k~)S�@���Nb=�$4���˕�!-M)d;}۶';M���]S-L���mU�\�{;�v�l�:m�;�����$�X�*Q��o��%a��<���u��*��3�(����l�ܫ �g:�K��3^�N� ������{S�T�} 28E!�!>e�^��
��y���}UP����"�n�L�B�� �<	��b�`E���7�mlhɰ��w��|S��%�u�ϒ��Ka���2�P�n���>mQ+�Vd��<d�vm��E�����0^4�b��)k�.jGd=҇VQ6���kg=�B�@J�z���?�h/�&x�l�am��� A_���Sa������e�"�ۨ��9��<كp�H��12�Qi�FJ�|����/"M�AGD�@~tv�VJ���b��d�Ȯ)�g	�H$C��x�Z"Q�U�D��E~��Ԡ�ܞ/��{勩!ČW~���ЕܜEx<�������	W��y�p���dg.������O�dF�%�6�����;v�P�:��3Wb��PL��3���r�	��_b�a�Yoѐ�|��%��hKgmL��6Cβ��Jra@�p���ОF�,X�]ڒD|1�û@ƺ��+>�@z�+ �tx�p��jB3�x���j��$^����F��u�mF�g<�ҍb�2��]ޟ9����`S*)�)�t��\�ە��	30u����`�)���ҝ��j��wa������G��r�4lG�ݤ�F�u\��:6:�����b��� ���>��Lk�u��'||�H�E�}���~���y��u�?�r���I�@)P*m=�?&!=�����إ(N�u��TnN@IHO߸[�wn.��3���u�6�0�^II�@����" �������+�{I��[�	��7s"��q-&U+��$tщ͑��i�a���!`��=(�s��1	+����Uܺd�j���߃�CgM@S��&�]��$L`�/ߤ�B!|3d���ᦰGH��&j4+�.1��L�A�H��Ać@�4	��ޒp�ó��u7?jO{�>.�k��Z�}��so�W֕��������7�L��#%��%��w��a�֞k�·tQ�d\���R�Q�g��d�~�6�a����cS
-�?%�"���,#n�|t�*��y�fK���<q�
�|���k]��߼ζMD잌��)��Z�Q�A�\�c�{e�8�V�S���WY2���	�##�^s��h1�}�`r<=3�|�K�Y��t�� aB@�!��7�z�.�,�{T�;��2â��Կ/'���%��\�� vi}*�1H
��n���N2o ~�z`������(E�{t�.~\t��������!Y�\6B��8H�c�uQ�8b7Y�> v4�r�8�&V��>�%B�W��ˠ�M�*¦~����`t�Z寕[2|C��,t��E=LD��$x���Ϝ|.�*%�ҭ�R��%֜�̏ߝz;�ҭ������/;�k�;���ڵ�����>+�]��ؽ��q,�֖Au��&�Ț�E�/4�3R[�����[P���G��&fV�!�|�L�Ny�I��;�@$�$� ~s
t��^[l#���z�vO�1���&q�Q���ks�]���N��"�������\���=�L<�����.����
�4�	N7T*=�rSi��cLq�M`c7��ЙlkV�|�LH4����XK#��j�Y+���b>;���X�:�F���#-Ac G%�����%��/M֩?�,��ӕ^�s���
��������Љ�bqN%"�u�w�;���=
]��׀{�\������ c*���B�58��бH�����Lmy�����O+��U��̃��(��$�H���IP�Dz�@]�2斈jCڳa	R�?�SS]���G'��{��8��0
+��X���Ϡ/��Sns��?Hf�d�sx*dM�"C��V�{mW*|�h��^�m:I*?_�4�+FڐN�p�>%*����|w���:�-�݇	����_�6J�k������];����[E�zi��)ȅ"����8�|�Oa���c4�l:��3Ն��U�E�$�E���ڰ 8�n�7�����.�z�4��ˇ�d��6��0��\�%#���$�L�d#�މ�%t��_@"������.4F�] ��H4昉0��ғ;GZ�L�_Ќ\��%(�Ɨ���c�N�.�j	�k�e�,���t4�������v����:^���6��ʸz]_^��ᱳ���N�N`=����x��계�N�	�8���� ���B�+NH)C�T���D�A�u�aZ:�O\WÌa8�x�{d#A�s�yx����[u��wX�}Й�>uN?���2D�Z��7� ��©��l�+a���B^�h�T�3��$�
mĽ�e ��Jz.�~u�o��V;㞸%�7��w�ϝDP�z#��N (g�t(ưf($�1YL
���X�������5D�G�bVװ��D��i5����܌ @1�V2���\Y���X�M��ʛ��E}T�з���Z��=\� P*�8�yT��B/��fnwhxd�1q�c�`t�qi�V�� �+!��P2�6E)d-�	)�Z�^}!k��m��=�c��Մ�~>�K�̐��6���@�>$���=���:hf�ĵ}�p�iQ��:Xg���1�c9-�(A�n�G7�x�;��x3u ��|o�q{2!é.�ʌB���
�S��U����
{�j�ֈ���W��0on��a[7B]ϹJ���IH�|K��y5yl$�p� �Х�wPK�NIvP*�/�̥N%���+F|�t�%2� +$��B�I�.ʴ���3����	>�������bҸ���nha\�Sx2*�4��?`"y5���,�5}�A���Eq���?a�ظ�V14�Nqw<�<�}i7�1��V�7�l~�!sq�b�1�Z�"G��э4�^�g����7���U%�]ė�K��7�g��0͠X�O�>��_��qc���07���6$��J�]}Ɔ�t���5Or�����0a�� opQ��_���d�n���l�J�51����������8�{`y���p?��� )S��d���1��\����&��ɮ|C�9y�
ń\���C����"�e)AR��*n�:ܹ�l�P�nO���O���_����yx?��Ɛ&�܋
Q:7�u���7�����A�9�I�_
g�L�I�����V�v]���j�~蔱�>QnS�
	��Q�d(�E�U���$^J���%�_�8�!�b�A}�x\_���'�h������;t�{	�w�czu
T�g}�LI�.�F�)��K��X?iҲC�KTW�J׍��,���vn���~��؀�S�����i{z�,���ˬ(z�{����I�Ǿ��T��Iu�?o�����b�a��X��WdTBň�n�9���}����ω�9� 3�����o����d�J� cMA�b��*�(s�L�
��16, �A���V�~t+	��b��	�������������	t<�a�c��X��V��
î��!�@/���3�\�^�&�,��ڼ�h�?*)L� �����S���T�Z�-E������`�Α��}X�R*IW�XL���:{x�3V���/�+�G�1U��?��$7ی�s���� �������Xrs��Y����嶦���I8��������>���4�$j�#i3�&���US�/ ���-�s`�W��`N>����ǹ���qb���b�f!=����H��x��GVT'W���q}�����ҞA��R����O��Q��� ͑Z���ڤ���o���S�{&����/�;; �?�+|���T��Ƿ�O�V�#|��B_����Ha�����2�W��ˮ'ޠ�,�b'�똇���k�:&��,�����9t���j�V�kq��`Jz5��#�u�p+�,繙�5e�2m�����R?�l�/m��*�	���r��E��x*�#H(\*?��iB��oO;��.����d��v`/�}���L���L��<���J�S��+�iZ�r��7e��LCz2+��6��C�e�ʻ�H�.�@	� ������Ģ�������?�6����&�h�&����	m�f�l��ZJ��V/��!%"�{���_�
�b�(��qJ;����M�5����Z��:2�u49y�}5^0��ߚ�-RҪ�O���Lz0CD B`��s>JS�i\96���Ե��(wf���^w��#(�Eu�.\���>Y�F#A�,�5�/��xi_��:�ː3������S����Q�H���l�����4���͉�[�G����8�M�f�29
�?���(-dXO.۫�W�\ ����L[�n�ӻ����#������Wc��s��~q��O�Q���0d?/�Y�b��Щs��S�t�tb���C����e6��(P��ZR�5uX�Q3?$6�Y00{�N09�U�bυ���u�Je��-�l���&da{X��CF�m�y�����A*9A8MKfUn��G�����)M\�l�)���v^&
�du´����W��<�����I6��Xh�������I�j���v7BՎ�g&�f�>�EI�)�I��x�. �l�TJ��~46���SǤV��;)�:�>�2]q�
�֏��S��ѹ��:���P�gjo.�ޘ.�������ֺj(.�8�9s�����^��y� �>A�S�?s���35� R`�%	�_����6�п%�R6��"'��!��v 0mK>��q�����)��wI�Q��W���M��ie�v��h�N�6��P�w�d%���T-qΟT�{�r�>a��@=�B1�y��b�w��/�v�IUZ��
0��Md.�>H1|?e�jb�oG�mC��Vu�b�VY��`�2
�0-��`�7�iֽn���Q��Ѷ�����D��t^uO�n@�&Y�U���I�Q	bJV]��!���j�y���{|������)@�̈́�S��� �nyK����{z�mm��ч�Sc�y��U��.+�P&��i��Тۼ�Fw�<�;�M��],k����c�p��q{�w<g��p2��TP�F^9Ц=]3�<N��g�|���_; �����ޘ�p�&�� !OT�	�R&�O��7�r��}?�6\��I`>s�K�LC��H("�2p��_���E����K���6���r��DHz݉���'�tMyC'd��C�a��%'Z߉s�H�Ğ�7 ��@ ���g�a����ӊ�+��Ǜ�.�ko��y��Zڂ���L!a/��<g����2qJ2=����j�A��)��V3/��Z�AÊ���d�_E��<�g�u�}�{x87����Wc���=��*�̓���V�|X���oT�#0I���%p�����D��V�{yV(����tj���T�e��U�po���]�_���^gOH��}&�D��}(4�T�ˊ�?�N�aZ�?����`��w�k���QZ%fb�9o�R�P�.9B��/��e���<�[
KwK����vX���T*�������kh�>���]K�8��w�~��hHY�Z�-?:Q�Q���:�V�Թ`g���4qy���U,\�m��s �|���.�7>���s��$�ѭ%�K���R�wo���j�O̥j|}�
�(aR�հ8Eݏ�_���\)�3]����!l��z����!w����uy3�ź��U��A@Tܸ���ux�b�V�p�,F	S��z��a�w��,>��>J�s)����p�t��ʭy��PL!�7�w�D�&��TX�Zj�����9�~>zn	�<��o�]&�ܞz{dTp#�H��0Vc�`��=���o�*��2a.�X�bZ��JS"`eɊ��}�<�u���ɔ�bk�Y��<,Da�*k�jV �3L�M)t~�,��PӴ���U�LW���ת�L�,�d�.Y%��S���^�� ��vl~ҁvՏ�Ϻ���!�7\���~Ge?�zRP�������:�5I[Vw��H�(�D:��eE̾J�̗�~��E�"���[���=���ךY����y��ym��Ыr���<��Bj׺���6���}5J�q���&V�eG7aJހ�b�D��5 1խ�W���򣌘A=�/�/i2�.׮��#Fˬ̓|C�-��>��)�&�ҹ��T����B`aC3�Q���_�#]η��]�=��� �\�S7Xf?E؇�d����[�k�SK����T��(�0��R�?j�����Ak �qB���*^#�T�j+%4 2��v�����h�y��:t;�D�G�W�P���zb�D��YQ�-�������  U�'��is�����5��\��٥80�1�X�� �'̃�F�k:M`���Ǡ_r�U��*n������v�����ڻ���2�1G������Q��#� ��Ӝ��K�A�<p�!�W��<�]%�gɏv�<�sE� =�W~l`�j\f7�6p|����S���c�Pp�����4���4|���z���
���Q<�{���9k�P+<Lh�p��P���a}i��z�:W��`����se]��!P�J��X�5����1>D���29���#��g�?\}A�$c�d=��R	o������w踷�db Aa�{����9�3�� y×~��m�c�P�Q���f�#Jgb9�Ǒ<|��J�L���G�n;��!Ք2>�qF��>
�"IA��amL)a���͘Vˢ�?W��E�!�J�٠|+�^g�Ti�M}ͮ����ã�ы�
�Xߛ������ʣ�f�S4�v֍��{c��:8�����<�����Ғ���(e�c�h9��z�a��
��g�b>�!��b`-�s�I���O�|����ޔ5\���t�'���ʪT�:�Fq�S�i���F�v>���`���z�������"1�qgb�q���l��+	h	������9��
q�ݾ���լg�o��R�~�,ug!����Ғ���!�����˶(~ �܁�l8 K��}����� n����G�:{���o�����g���p7��L#�2��sE4d�/-&u����U�U�x��Y¨S���
���nR���Wp�꧈�;��@�����	&^[��<��l����浣�^�{zs�a��-����= 7Մ�	��Zy���A`|��J��i�-l�����~}����������2�Ų�㦟�V�󗝮9�'B���R��}�t��\9{�E/��@���<_=�@�SS|���-�ԏ�X�\�^L�%%��{/as�"l�8('u�=	��#�C7�Oh�����+Gc<n�'�Z���e����e�er��3��a��wKa �����%n0@ O��L���^9����Z�XU�X�wBS`��;�F�a*��qtO����/ߌ"d`��a�����2�5R���@��g�G�Q@N\���CN��pr��{)UP�^׉�̢{��8�l�u�X?5eR��BU~2����q��;�gj�B7��бx�EF�s��H������o[�Z�%t.�����&�Ҭ�P���juG�ZuY���S��q�\�f���!�q�*�s|��%֭$��:�Q-,����|�4�-��5�����,����Zٖ�SᲰ4�����S�l5�9�	j�2hc>�����
�����7#B���!����"����X��N�[�S�jWOQ��3{*�X�p�/B��`��l��-���c!�u;N?�I�k���
����{7�s����e3�ͮ�-0d��4$d:R)��zX\�5n�0�o�c��`9��l�4��4� :��9+��� 8����s#e��/b#!.��L��X�Ґ�! ><�_=����-���>�^Ҍ�K��,H�^��U1	�]̯ #�ΈDԇS�g�BҪ��lA77�[������;��k�Ox�<A�_����%�ksB��mU������]��#��w��F�7p���J,'8(C�>�!A�̧�/��	>��ם����.o>�ӯG��7l̰t��`Ӫ�Cd�����[����z��6+��נa��j��]<lFD�uL00�^+*���e��Cx	@�K�B��؎ګ5��=�cR1�������T8���1_,�d���gM)�*��4��X>�E~�)f�7J�`r0Z��R�?b.sG�7�H��0�'ʏ�6z�tO�#x����\ ��\��FRa3 V�E-/4|�x��A?K���ym�i:�Xap���K���ʗaK��B�qT��a&�tw2�~݌��1�"�>
�o�Ŋ�mF����+��7xm��|l�{��S,��܈3�	~�A�0�GLa��tE�@�»ւ�_�s8�|	h�"'��IdM��L�ބ�WM�]����[��)�޼>sm�Ǭ�R-��P�tܫ���m����C����8�+I1K�O�e��Y���cFO�sS�.��i���5��8�p0��c	�M�2��:sl���$��)��F9�&�"����;N|�\��q��\����n�ҭ�`���q��~�%��
��Uo�%�?#p� I��܄g�1�C���G���L�?ES��@����/T�\�_�i�E� ���M�m-��W ���5��-�wfzgMH]ٜ�g��Y�8����5X�&i����hR�E�$���
+���4S�+�{� g����7�do�$s���)m��	�W��K�N���t9��]�FR��t���6�R���K]���2<+^>�VZnx4��N%!��|��n��a��q	P���t%omd�����pgf��m��`��Ky�~�i��ʘ2VɰMI�յ[\�ͼ�����X�:��*夡���o�zV]�/ж�B���\��/�@�Ҙcet�F,D2�t.?�~R:�M�����s�Ų�Ue��Ef��vc��JA߮9i��c+֢s�5R��-^������)�:\�Q���#�h(���J�4��&����U��y����1�v�.��{Z���
��j�Y<y��c�s�.K��ޠ���a}^0<������������[��� �`}u[v�v�+c��M����#�jm7(-��lM�D�T��W�zX�,�yO���f��'w+�iw��҂��ܗ8wi����sG�Nb��!�,?b��T�{rn�<����d�a�Sፂ�;�>���f���U��6:������	z'�6�`���,��H����a?�S�þ�YU1>B�I��!� �N�g��ؤ�Ӳ�F�]����|J���q����``��c���`��&� 	�}=n�U�� 
u��Kh9?d4���"uu"I�3�}H�����y���%����������1�Si�.d�/�}��}(��*�|i�洷��9O@�$�h����
�������|.�b��@�h|=,������5W�'2�K0��E���־X�|e@}���E]?j�~>�rB��z��+S��I�#�M}��T;�nE��0+".F���LUQ��+e�~ih>��\�5��#e�LsU��7�Lf%���A�x5ux�����ֵ7ǅ'�4��� *ii����Y�%F��ߍuڪ��7m��(�}�Ǥ�2��ݤ��vWPx�`�g�a٫4!Zj:����l�"aQ��]`�H��U F���`D<��X��n�B0��5�G>ߎ��d��6m*���<u{�VF��N��4f#���P<u�Z�4�zo��vhNc�
��<O��ʪ�d��<�f�c��ADԊIChc9y�� uԖ	+�����g΀4�R��۝h�{���>W3�c9&|u��1x�1U������jI���IκDyY�x�`:�آ�GV6x�¸K�A�������F�d��8�H�zw�)<awa�L�����l���{�G�[�����nK#vV����H��O��Id��{����G�!$��]f�6�_�����A�eF��%QYʶ0��3B��$�^�,5�ċ,��l�ت�s �h9C������x/����ȁҳd�G��JK(n��uO։(���|搏�U֕������k��}2Z��TF������,Z�*Js��w�-.`z�;��.�@�̰���X~F"��4�[6�o][���[�￳�G=��`hy`nxRyň]f`9�Cc��xg���n����͵�V��4�O��=�u5;u�4"����ǥ%�^\�׎�Ȍ1�Io��X)�mb̋�=<I[>O�248��y����NA�V��9]Uن0<dޤ��j�aX����pp}!G[%P���y��6�2~�~�e><-�%�2��I;4c��gv���5�=`_)�W�m�w=�=�<�s�+��)e��GBx�.y�+�8�������� '��wU�O(���>ohc�T?{-�	�g+(T{����eA'7��6}��6���2���`]#R��c��1D�cB=���	��B����fk<3ǁ�5
��.�}�?LM6�X؎eL�帬��Wg�NZDq��!Y΍@�7l}� BW��� ՞�����RFƝ�X���ؙk�,�����ɨ��[�X�����e�U�kϐ����t�����'�������ΘZ+J� A�� ]�e&I���.P	:��uGltq���0�$�M��8�2�$����N,+��p��cԒޓ��S���G���5�B� �G�pޤ	�5cK�1��_d�V-Z#>�I���ʹ>��s) s9>�nGlē����oL3>.���:>|[f���X��B0�X�̖@ �ad��'�z�0X�����'m��G �xL�*!~@?��������_IHG�$��ܒ�2�F8�a� �G���_��QR��������MI����-���5ql�D�X��e�˯��! ��}k&$��07�h<��������is���a��0F,���� �舥<�T���u�tė"|>�a��Y[�.��v��ҧ1iup"��a+�i�$��n�2h#Vp��Qa�����A{�.g�uնD��
!_=���p�	��L��{'#4��`�Ÿ�9!sU⋁
���M�G-I����M/:�
o����*�8e ��5��a���u����9}���	�4r[���{�s�����	i]���/�ˮ���|���6����#����ۺ�$E��f�M�rB�����͹�աgέ$\�,@"�-�@�W�3�'G d�ƒ�D����T
?���L��9��
��̛c1�).�C��/n�D+�_��97��U} �@���I��kQQ�){�j�kVʶ�%��s�3d7 �2ݵ��[�Gݙ���4eh�H��ˆP���Ǆ���W�-7}���_���5��H4���4�c�H:0Pb{o�.�z`�ig{�s�Xn�-H���-@�|��K��bb8,,pUn���Ycy��=d��k�4�׳�m�,C�?jVZ����N��Y�;�D8@f5�)����T5����\�����ZtS4�1�}Ӆ
�%�͝����
KV��)�
�'4<�	>�Ķ3�ғ�'m<N�`h6Ú����ӈX�	o� �WEn���QBP���5�"�����x��:>bⰣ��D�_�Ty�ɶ���
s��L�S1E�À���^��wY��m~v�#[�r��5 3	k�`4�3���h�.��]�%s�
��׉P���9d^�֘�z?3�'�8����@��X]�l��v��1I�6�m�.9EQ�/^���F>B�PZ�j��������cDg�}H�xWý�-�h�h��X�4���J�4�;/�Nz��p�p�j1E��A���}�%<��M�dzp2I$?���� \Y�a!oSsZ�*�8�u���+�T*q��5{.&����笅�E�@c��VK������ �"���!��u��F��x7Ȥ��eǸ-o��s4c�k{�pP��i�k�eX����l���e� oi��|�O��A(��#v�!�d���iIc/U�&�y��X��3<��W?)�B���� 1�IMkpElU�Z���
�[����0Zz����Oq�%�A�<� �����J���������q?Ii5��N�$^�k�й���.Stx��S��գt��a�k�j����iNX�0WVǗ�	���]ҟn�q>浤}Wڢ�����V�Ϫ.>fv���ä
F)~�X/�[>�1=d�K�jw�����튭5ez�mѷ#ֳx�-a�Cʋ�ܢ�5(��̧�W�W"B4"���}xVr֟		]:Z�R;`	n����2��W�%��+hq��$Ok �̈́g�/�;������F��{	MQ��Zk�N��k.[�M�g~Ͼ#�ք���3��X$��#v��J�ܞzm�)�M�k6O��a�
���5�!�y���맣�(댝�0Gsp�ٷ*Z���I�5w����-Q#���pΡZ�����x���<�ۯ�¶��-��N��*�R������G���bzH-����huRX:����|P���*��/�04#����2H�yl���g+�V�����=��b`���0eѣu4P��m�8���qo��N�x�����Ĭ�ޅ�i�������9�C�)�0���6wY�G����j=ü`�|�}�MO;s.#��Y-iT�NUǶ������?P�ems�k��`�{���MD�6�F�=�ްe��K-+'�������L@^��������t��l�P֌���H�<��L���"�i�١POi֐����}�Q�)�4/m3P�����`�9!X��iiQ`�[
�g�O,�|���j.��0�������'Ň�ɟ{	D^w�����δ�G��^�����);��\l#��T��I�XU.	�LfHU�iGc�} ���1�揟W�"F�{`xY��oo�J��2���p�V� �]kOrD���lj5�]rtV����t�M-tx�E�,���zy�����V+Y�ʧ-\�!�+��g^�J}���}���������ɠ¥_��lN'Ќ��Z�o�����OϑН��T�g�����}�)n��;m�@�~}�	�7p�g�j�i�� �����A��������y99([f��bw���:��Ed���Ҥ��#t����o�`��l0�5� �ؓQ!����%�{�K��ܕ���������R�� �*	�)$+J��ͲFٴR`0ņf>'Gm���[�&u��z+���V�@���n���{^�N��G�
��#�:����R'���Z��,r�+��=w)�@��kJ���K3�i�$�-�/ђ�t�Y������u��K��Ǽ�(1n=?�ofU���jn)/d8A~.��k�gF"��C�,�0�`y�|wp�W���8�r�;�E�:9�ŏ����G�]�} \}�]�{R����k���߹I��|�TQ`0��O�+vS�R�1��Us�d�[�E�_rw����~�R]. v{@{b�}�VC���6��'l�$6��6�ɍ��δ���(!�^�5H�R�e~�[�<XW��a�tN]S�|Q?�5�*�2^�Z�(]o��>dV�@����J!�}���A�����3y�/�/��.x��P�w�����>���.�3���X^P�\�Tݤ$6���W� J��G�.��:e��<�t�Q���ι7^�����n��|�bSh���~#�Ն�5�vp����BY����q)���,��C������R����l�3��)	�dq����B�L��`"{^._��.&�,P����t^W�'��p��H����w0�������N�L�g�չV�z,@��Kob�k�!4,?�@�΃x-&�\5=X�m*՜���hbb��ʲT4�F<9-���T}��{�8
)$�B^�"4g}]y��� N�`���j�DT��bU+��cο	ߓ:W�ܲ�v�W���w��Z'���<C��I��w*A�V~GY�ɬ2���_�m�Ǹ���l#�h��~���gjsQ5��>`
ic��dJ��]�Uv�؈VQ��]�-�J�C��Ϥ�)�$�<?R�╌D�םu7�%m|�U�U�d�+\xyH���*�j2�3�e�\�ܛ\!H@ETTQ��?H��ׄ0_�(<�V����0�1S�~<�1rmz������)甝���s���TǨ`�@�p�Zu5��9��?���4�RD�<�@��Rfr��%�`wC�X�a�m��}>�'Ե�.�jʢl���ޜ��_��:�8o��Č�tk��W�mw=���4��9�G�~ڍ�v@m,5�b�T�BI,����N ���9����J<>�8M+c_�V��:�ڒ�~�_D��Mp�J�ds`��)p�=|˓�f1���޾W��T��t�{�v:���� �09�E�6��$��#s�O�t@I���]�C4W;N?j8�7�Y�����&Y�j>s�� y��P�	�#� +�zps�2������(Y�O0��1���L�k��i�N�ᬀS9��h�(�����샰��#�/��K	K�gI
ăx���D��ٔH셗�Ƕe'-6m��--u���z�np�ѕ��Z
>�*����Km��#�PR�����Ͻ��������C8�צV��D, ��J;>�;ѸY�U����G���F��O��@�M�m�.�K ���$>(c#+Nx�e	o�CX��}���2v�Yu�,K�_@R�� ���׎LD�D�Q(��rWr�ܯ�n�#��"k��!O:�ŪM�����o���<�,z�Ͳ���p� ���vW:�H��o�Hރ&N�qc��e��밪U�쇃��Y
&�O�$R$�&�k�)W��l\ʿ�`QG�31��I4FA�Bu�B��|y�H��+�h�ё��Ąu�S����L
#mΗ��
��bh�J>��n�,->V��Y������"�A�S�,��]��6FF���ɋ*4�4��3�L�p&|�Tb��ES��(3��_�!��o�,K���aP�^H�i��o�.�H����,���8�hb|��X��J}�
�����]�,�5���CA�t2��mt�P"Z,��odT�laG��а}���C	i��Q;}�^�+��(�?Ē�삜̉�U�Oˋ4H[��f���x� 	s�K���1�H+�lfM�&�`�N��$�ކ	�C�>D��5����Cu���32�ǡ��`LY���!�m�Y:}A�Hʚ���=FZR�-���-�[��^�p�����/$����_���hH�˞T��`#��
*�$�@�0�z ����a��5���6T߇�6]�j� ��we�Ϻ/p�um3�|6F��q���/+[�L���s�a{y�n�����ȥ�ݝ@)26|��-$����X'z����B��i�-ÿ���
TC���{7���X+����jnZ�G��q,7�r�%�@���#��+I��CL~/��؎�y�墉$�a����&�!4�x�#���]3%km;��0�E6|/�(-�s��z�l�{��ȭ��,a�шV���u�u��,�Ȣ���'�l8rv�}"zIV��@�JMLYl �n�'�f�a��x�� ����c߲�jVi���#�[<6��-���[ Z�,�_0�7M֥�0���a	�T�Ʌ�7�#���[/^��Nxσb�Vx��ς�uK��(�����YҧU�lh�6�U<7FP>2���z����� ���n�W�jq/H��=M��t��q���l���,$�ި�p���iJ����c ����Fe
���Т�H���͋�)-c3J*�S��\�i���PP{�[>ӣ!���}���l���A׀�S>��'��	��>���`!9�.���;��e�x��Fb����mq	�4QF�����Z}K/��w��2��<���Ǯ2X�2��k��@$� 6��O6>���%��U���P�
0�;�i�vQ�T��N�A�c]a�2�����/��ZB6V��b�UO3@�J/ ���V1B4.t����4K{d7���R�G��y�)$�Q�����u�\�Ѕ8�t=�{�כs�ƿa��Y8���Yu���������C��l�vĘN�0�F�����z ��̮sw���ߓ0+�-���&�ǲgo2u�Q!�:����a��g���}Y��F��'�BĦm.�[��ƕ��Z<}��?��-���yF��jK-�U" G,bj�h!o��qL(
�����"ֱ.�x]��{�IΛ��C%�ySxh��(��`���#�K�d��ȹ�;A�O���a>��[�o�Rn4�w;B�>���Z�W
���gyF�]u����{$}ڹx4n73
^e�T쐓���1[���JXY�g��OQ^+ڬC@$�ڞa�b�O�	�ܠEa�1&��P�w!��q%����sW�G]�����ޚ�'R�\VS�~܌I�a���6Я��×��a��}�A"�|���Euw��2{�p!H0�B�Vd3.S�o CUy&��+��z���_9�G��i��WC�%�]]����[�5��I����X�\�'w��6i��$33^��&Gg�N�"�l<�Xt#��ޢX2X�����V���Pjr�W���-�2.�j�$�	8$�@�ih�2y�FӲ�Mˇ���}X[��m=����+�?ႛ*׻�a�|��;�4҉�0�N�%� L=N����I��j[�4x5+�U�b+�׃o"P醀��	��+!γ���8����:�MYݫ $�`�`��	��H�#cR9�e��h����(�D�}��]+���Dt2HrV��y[ن?a$%��S���`l~BP��1w���"T���.����+P�Q�
.(=���h�\����<��۶����O�tR�Q���t�f]zpt9���q��3?^?������
���CD~iJ&48z�ƭzҖgK����&1o�r���}�����	2���?*�Cdl�yФ�HK����o_.�	컮�4�؏J�Y�&�?U1������i|H.������"M~10p�t:UT#��?�]�c��i�6��qbÍ��T7.����<��	c�{/[�Mi�d?��J����u^i�r��+��I��
�$ۺ${Q��/���Ra�F��7<�l.uc64����%���@ht��#ϙ�%�՜�Crͱ��;�ЪG�l?�<�E�Nc%u8�<x�Ϝ<�`�O/L�=�����xX&eT�>��D-�H��D`�t��͆18OP!h�$D�&�F8��d��pJ�
+��eO縑��g���=H{f�
g�A;�*�H���L���9�lAx��Ƹ�#��?'��̼{
�ю��C�
���T��6�"�X���Uf>��\�����aYӱM� ���/�ֈ=jn:Ģ�~#S��3iVjڛm������W�@O���K�Oj!��~9~9�9���^��w$�B<}i��]�91J��T��T(áv����PaX��,#��x�,.!��(��t�}�udt�V� Ji�t�u���֊`P�6]V ��)�bqEob(�)0>�H���W)��}%���3��+�F���=���A:%�2��2��q�楛[��S:!#mC��^lN�XN�~��ORjc�:C�D���Zxe�= �%�"�p�Ê�Z`}�׼:��{e��\��Y,l�@��z�hjMm�Q�d>�Ш�6��q��1����.c�1�z�-��(-Z)Η�y��2��_oa�:����T��q0�xq���I2m�QT�N
���<��8&�9,��2K��Dg�Ƞ�%~>47�Oi����xu<�p�����>6��"�O�|�q�����@�劬/��)���;g�����c� 츩O��4����mG"'2{r�1x��bl>>@s����f�����t�YB[״��/.���X�`�H|� �������O�����h%����GٕR��2=CA0�p�amuN���ןZ��ľ��4Z
 �u�̛�;K^�.����18,*O��thi�쒍�Ĩ���m	�ߜ�xj��.Y��Y��-*��^��8��[���S;��h!���%�k�������遉�+is�a_�U\�G�<;��[�C+r.�����f*�
����4�,�j��������urk�Z��sA�?ͤu�S�6u��Ȧ���\�ԲJ\ۖ>�Md<���0�s�ɧbB�o��mEX1��QC�����D���ւgѢFqw�>ƺ�%�Z&p�wOߠ���f��S��~$j;p�9Au��|/!�]o��H�e��w�z���c�$��<s���,(�)	�ZY+-�r�֗������4S�ԝN����ICz�;W���uƿ$?�`xW�������݊�8���-Ku�22y�t��r�F��G&�q�G��&w	k���s��վ�>#%�-DN�6�T������C�����RKsS6�!jc��6����Y��]`��.����у�8;��'�Y\CB�m0hA��-
3Bj�s(�{o��d����<����9��$��ZpgΎ���0�]o����|�Eh���Vq`RQ�ت��R�[�!3hsl� �/�F��T��
������2��@���:�7b������l�cFI��~m���5n(��lL�r�N�&�i���-�m�b�"���_7���!���*���W\��E|V��]Z]U�`��x&z���c�P�g��ܮx_b��}�k�ghf ��5?u�r-ˎOZ�f
����b��)��|K��B���#�$�ئ\��,^l?�x��R�S8U%*�wݪ �/��y�6�w�-���M�!&�A�"8���%���f��o+$��O�Q�q�V�,	d)�8�c��%�n��G����Gu	��P�h��y���S��l����%z��<�h*v}�[�k�0�	V�۶�cV��@s*AEcQ�<Y�6�I�b�<q��f0(�T+�ȯ�<�?fZ_�e;�y|j�i�h���W+k�=A��r_W���'��ˍ�{��آg�*_��I�3�V��{�;cb(x�-d����V�MaBz����*1��qB�x�0)����� ����sd4����2�����ɣe�#�y�R��W�l����m6�V<�����}w�UݞE���G�Ki|���!��E�%�xz��(K���_�5" ����攱:O9�D�c��E�W��ԃގ���`s�J�pE�qdk���E�@�:h��Dj兤��zqW���\-�a��E����4�뒐����r��2j� �P���_�����d=�1�y�<R�����@ȍD	U�bY���i�w+�P�R��L]��(��h+m�t��wڇՐ��a��W$�چ3��������Id��#���9��A������2X�c}A%?�<�P����M0X	Ν��ϊ�"�Ǘ��r�5Vb�C*P�jb��tG6y`i�ddsn&�n^(�r%��/\�tI���4�� �{B���5�Y��J��YB�L+�;wT��u��?�:�M�7�1���8��Z �-n�Y ۱�)^!a�S?r5� �&	G�.
'A��Vh�wgS^��+��gL6�+6���pI��G�b�������x�%�v�\�#��	�b3汝�p��VuƇj,0�T&<na����6�W3,����R��ņ^����T]x�q�)`��ّf��H"ŌH����� Y�ew�.�s7Vh:<a
�ݸ�P�������=2��*x�])�]�C�@Qn��	^����oA)����6P�` 2���;Y�nM��İIYN�\C}E&�UV�h������r��qOԛ�M�H`�E��<ڳ5���{��V/)�e��>,���\ FɈ]�:��'ҟQ<t�͑�:<����
ܩY�\
u��Oò�K㢳�m[�ͣ0sF3�����Y�4N�|W�|0d
]��D���9N�n�������>��
��`b�m�P�p]OYr����tx�LA���B�wƒ�ɂ��lHm�^ǋ���ח� /8��ؘ�w�7�=[���P�f[LjI�:a�'��2��m�o�k��3(���yt?p�L�������1�#?�݉��0t/�K�+.��q�l��%X:#@�J;�_���ݱ��X�[N�K:օ�hŅY�pCo�"aT�j0x�X$��	fA�
�����J�t�6���D�-޺�}��\^4E�q�,�Ϧ�<���t��߿_S�0�jQ&T��t����w�ZL�ҟΊr#L�n������Ϫl�^� �'llz@4-6C��	�v҇0�q0����y%2��/i�9��� M)�a�y=�3ʶ�.	46��c�3}���S,��ix�3"+[�l
O�3/���������^A�)o���d&���=MZ��?��/�d��2���#Qr���)�	�����Ze��X~<3iEư��4��n�s0��ʨ�ﴎ�R>�}����`du���M�T�J'��2��]4<��� �����
��ʸgP�O���^��Vۻ?�o�w�;�q���?�	F|�����n4l��02
�N�Tr%�v>��x�RTp�T~ ��YR��@&�Þ�c�d�d�Y�m����L������l�Ԉ�,���	��Cu�Lgw�H��,Vuj����\�0�[Y)�mWɂ�q1����	h�!6W��`$���f�\f��w{s �+��_
����d��̫�]�����ze�����C�$���T?[�}��7a��b��~��0��Z�X��Zg6/K�g~/�����K�
fޒ�ni����f���4����F�ir���/�5���@zt��G���-F��	��cG\��~���]9�O���-S��X������t���ⰴ��JtrO%*z���G���=xGx$c��$C����zE{�Q��$�n(u�H�W4t�k��R�d�J=DZ@	�]��a�,��GE��ZU���ݩ����a���M?sW�;�y{��7d<H'r� �fg���[h`�]�t�<�l��a��j�N��f�J\J��%MOމ�	�]����(��	���tWֿĄ��*h��ts��K��眘�y��a���,�]�Bۂ��� 2g�!$�Z��2��;�<�t%.!3�1����j�h�i(&RE�l8���LET ��ƀP[;sr1���}#vG M���^�۞���f�S�]�}�i����k`'�9'�l�W�3�y��������[�����7u��<�Tq��A��6A� P�j�O��Ѷ�+�UPz��q՚�����;$=��Ky�W�s��gr���G�J�M�4'7�!Zk�MA
���1暋���.�Y�9�wq�_-9R����#p+cu�ZK��p��c"Ȩ5�+
�.Q}�C��3,g�J�����P	ڢ�u�X�e[��pn��w���Td���@�ܩzv�	���N�2NI&J��$��\�z��Ѐ֨j?^gX��X�z!H4Q^~����
�fe��m���O�L'���%�C[E�b�9�i�v�`%���U��j%I�u�ݓ$�)�����OB�ꁠ��b���&9U �	�L�%qY���X��H�7Э�ǅ� P-M��nhRϯ5���B�Z�GP)Q����S��=�2�coA�^�o�)�ȷ�*i/���z96�'�J�*��Y<P��"�*᫷^�������[I2������޹+-��)6�����b<}C�Ľ�4��.���/��w��̸v�HF./�m'C6��(��l���,�Iݰ\r$HQ(�}�u��d�v?Z+��JT����r��o+�T�9ɘ>�ی��}K7� ���Q�倹�>��S9}���3�ݐ]�~hm��[�,G����{�u��4!������8�}�e����]$\3�t�9�:i�Q%2�`F�Ky�����zA�v�w����e��U�u�	���(`aI���2� �$)�M^� ��'C\��ߌ/�1԰�z������iX���-O6L�+���i*׎�(|�+Psm:VX_%�Vb�x�i䏩���J	L��G���0�4�f��~1$��o�Md]��Y٘�	'U��O�����\��-�RI�7Õ�d�,DL���s�����^Q��B��cj�@�M��S�߻F5cF&,�G-�B
r+�K�(���Q-��ň{e�:�Y����`�`���~��l!-tX��$6��G��wE��4�*�v��y�
6��$�AՕC�n���L�����I3�g;0��׈�^��s�Gy��ޮ[h18�2Uu���[Z�����<�]�������wcL)lTWf�#�@l�YVҽ��a��|�°E�$U�N�(���ZK�����e��b_��?~WO2s�W�Q^�ς�d6q��V��{	d�p﾿�/�<��__���W�����.Ӊ�d�T�Hy����g��b���d��r���+��� ��TW�K������3��a� #Xl�AҤ�cGSGx��;�3 �Vf���5]�0�џY21<d�PT��x���:. ��)J���zaw(kA!�F��f ]S�Y�v�̭���UG��	2�g�rf��bm$�u�����8�mTa�H%v�{��O
F�MCm��V�Vy%��N�͇`Xn �GEGJ�5TM��C�]�!,��Q��C�'{��W��_�%�K|5�SgQٕ#��]ߊ��F���?m���'��H��WaeI�Gę��;�c��tRg���d9�T�k���eNVYR�����FWL ﷾Ζ�p�ش��-D'�)XjA'j%�%��f�ų����?}IM�--t�5#H�qcJ���Tţx����	X{�`�27$�i�y�n��F���r?�,`,n�}?��S�tƁ��0q#�L$DǯkE-/$�N��t�
Ӈj 5��q�(+<��w��!��0�Ǳ�J1Jm5_L����{���J��8i||��S��@�;;��6uL�m�n�pO�m��	Y.�r19d��O�K}+�����vg��g�g�t�[x�VJ��ԳP���0�L'ϧ�]�a�`T�����~\l�Q�&�q�4x�*�m �j <����ӑ�!��#�^���=E#���f:�z?fMl��������n����d�i�VHh� 7�� �R_O��h��B�-��qd����ɢ���ޓ�P{��V�������vV��	���;a�:#_��C�K�
���k��+��s�¡rG�r�\u�0��;-B��;����\���-|�H�a�t���U��4&硨��ѽ �>v_�n�[��u��v���J.���)�\�.*�R��U7��(Z�m�ʀ^�,�^����� ���h��D�/���j��6�U(��I5Ѫ1}��
�L0��@U�����/�D�~�.N�b]�>O^��Q�i��3��Lr��M]~��
�i�(��OX���@~���g��"j��b繸����r,�@�o�&�)�p�J]�0�@s{Yx�!�֪fI��Ey�k�_4mI���@z5?�.=d =��MU��D��0���Q��[N0Ҡ��t�f?�}������\�Xx#���c�X�;�%q{�*�d���;G�3��W���70CNuCc~�M�A͓�FsEtΕ��a`;[������a�?�Kx��Z���\�R\����;�5��}�0�#����Ȇ]53'm�<0����f�y&l��6�M�OHt�C�����)��@դ�M�<�]{����0'��B��� @��=�Q��$��N.s:�=' _!�/�2@Ry�7_,��v=(�L����Q�	G�Uo��z�@�䃎���>�����+@�1����R�G$�wVfT˲:�m�'��z���tQ�s��P�g�:��� ��R�9>�E�ev.���HK��c��9���U{���E�{���bwf&{((��E'A�Zq���jƖ�O3�U�(�DJ4�R:(��� �9���ri�.����%���@ы���w�s^��M�rm��LM6Fh`�9�	qq�7As���^hyx5tk7جIA����x̧�HOh�C��Kk��x�߀���hnǒ��W-j�ԁ�-I����?���jx)���Ͼ2�;l��3�	AcgA�D�g8�LFi�nQ���E�H�	JX���4����Y��^w}�����Jr�-�Z��I�#�e1ч�p&���_�V��ܼ�r΁
��I��)��$�d~�U>o�����Q[�J�G6��c?��7X���HB6ہyW)��W��?i5�J��vS��xd��57 ^�+'M�R,AE�����t�$K
�tx��} ��!HiH�7o�L��Ґ�U� j�Џ�z"X��=O :$@�f�Q߹����D,�v���fe?+M d�������0�a�rꨉM%l�4X2�����
^��YU�(�Cf��_��d3Z�Q�>�����ƐTg��9��?3��U%Ţ��,�����J#����v��\?�0l�p�4_����#��?��m�r���	ј�8Ϻ����.���$C�tPC�����@UP�����I��n���̩!�ߞ
���FM[�`� L7���у�D��K����Z��I�2	�������O�����6`��}�i\s&��t�o~ޞ�8+��:����*I��Z$�O��I)�f3����h�7��������3��N�,��b�iU!���۝"ZȌ�/�O_Pw[>^I��aZ�����PoN�HY�)�߇Zx<ac���q�9}%U�輟%�n��5�pr�g5�Qmu�(��'���%FAl�T� i��3��j�an&�d�����K*�������ƾ�*�!��z)�c}���º<7��ỳ:� �&:���z��2��϶ކ�$�￤\��2�E���y��U��,�3��rgpXȡ|*l��%Ul�z��٬�/C�pA�p����<枇��j��q��v�z=%E3�Z�kE; ��I��\Nb�h�F i��#P�ݫ��c$�>_*�����2��,R�T�@���J�����hD�k^����ةJ"�/��*:���q��[`�ے�]�=���[s2�U�u�Ԭ�[~ȵ�ob�������}���7������ܷ\���e�zҚ:�nKq1N/�T�3�W��W�ʾn��+M������4�
��!ZW�VA6�f� =���\4�s��I����E�@�Ѓʸ����􌜾��O<�NVSl-%c�O�1�z��0�l�G:�b�t���pr,���|By�Jtgeq^���4�[�����~{�\����T{��9�h�҃I�Ci�pA�̻���$7[���bw�Rj������
��Q.DLZ^3/f<�oKeF��?�R���QR3�z���l��+����(1@��h��~�*�W��������{pf�v�I ���;1� �������Jp^�N����0�����&j��dVմ�E���ސF�Ʈ1
(���#�}P1����3!�Pj�3���-�8�
�s=bI8[keZk�#�@ʧ�a�Y
�Yy�O�s��G���׭�ă���#;�E���M��+{G�c�[��2~�;�{T��F��&�1s)�E@#����}ޓ���2ŏ�T�J�q��hy���>�Z��ϑ��	!���nur2j��ED�� Z�;��5���[6k"�(97~�C }h�`���!u��x��$7
%�����٧T��	E^�L�W�����.ٍV��y^���c(_`��++������x��z���n��lr3�YElWag^���F�]J�Z-e�F���Q�=�s��ز5��	/����Sh~��
m�Қ�-�9LR5�;���G�������?�.����3�g8o�A�iI�K��}��:Q���`12i��ep�C�!XS�>�ep�� [�,߶�Ė�H{$}.�Ku����{AUӍR�)�OQ�������Vr*��S���=uJ�	�as�2������ڍ���}��P��b��1�2�&�F�GF/�m擏��������
H=�0�iZ�����ۢ"�[,7,��.�kPV�T������>�Z��UB�s��ve���
&2%{��n����R�_�$�_�e���w�z�����JQ=uI�!��:�J�s�è^����V7�h�i�T��.JJ�Љ��=\w��B�i�쀨" �a_���]̢n�'R�������&Mc�h�_�)�q�qMդ���2�s��o(�"�Z��%��=ɞMO����g��S��hC�L�ca+}xiH��w����	��N� 	u �$��V��!��Mn�EF_���4T�54�j<A?�o�M����ł�u�b����D�C$�O���ˡhJ�/�se_���PjU���������i�~�����q�W=;&�AW?�X��@���Q�0���:�P܋9Y��/0�6�v�+��l�D���J��P�~�MK��I�hG0��1�G$�?�[U�_6�����lP_n�Cko��^�I�6��ƴ~�oR���&�G��	�p^k�n�4n��^I��_2Wp��1�R��
l5u���ڮ�KW��̚^�Ưm������x_AuR�J�7��/�]�	<9��C����Y�4fw�`�����u;y�5�pcٝ"Ŵ&�����G������p(����� ��A�Hq���Da/br$�(^��v�$��FbG�#����.W�Z��ط�㉂z��u�+���WM�J�0�2(G�(�/R��ͤ�9? �x�B%F��_y�\��U&U��̟�/�MB���m�H���T)25L;0ZRϰ��U�b�6�g�2��Id:���Z�X���k�̅T{=�v���qp?d��
�%�����%a0V�@��<k":�����x��Y�#�����E@wk�oݗ�@��������jxIЃO��������,+��-��tm�g�֜��5]	�t�??��(jIO�)= E8M���e�n
�{s<��XԶ.�³�$#�EԽW�(N�5�!B��\�t��HvB�X*hy�c��G�e��o�@2��ģY(����j���.�uV�_Vj1��mV�\i����w¥�ܠ�qƳB�s?#�E3rr��o�3n��r����: ��d��h�v1v\�菥7������iLM�6�D�$�3�5�k}ad0::�X��:�ؼuv3�+��~?���q �o&�W{vz�0��5�d[���E��5�8�W�^�)�V��z�x�r�܃/-�_��k˧˱�Bd�g���&|@ߪޮ�Խ5�΀���ʂ�N�����=�����kCS�k�c�k@��֗kW�ݨXBc�<�$\0��nF�q>u��!p���*�V�
n��M/�;�yW�2�Y?1�����ך�\�~7������&?�:��t�l��'u����?Җ��T����#��������NHyc�_:1XM�B�-ހ�#>u��T�-��>uT9T�y34/"`P:��o�h��y�fw�+M���:F��d^R5�$����5�E���Q�n��cKJ�u���������)�����S�Y�EB6�0B�$�����Ϗ�w��؝GƗqa�۹M�Z�q�c��� ����pya]i�aH\i�Ӌ���)���H��^��t^5�v��rp^��$�k�e�(�xWW��/bA�s����_�:��e���U8��b���Z����:�����zD��x]���Y��87�+|�wN�qa�LI��Cړ��+hf��+�Ġh�69���
��P;kSj�(凙�ȉ��HB�s�ftƼDSO�����=Fc���)3��K����N�}B����{�`}[A>@�ʞ��%�Cl��/�>��9�����33
T2��}Ԛ�4~�w�"T)d�ê/g��~U��TlI�z���z\)pg��u���XJ���	Sq��o� xI��T���.+z�%��1vhѻZ���r�s����/N�s�u��#3?t���s���"o��p�4�|&'5+X㉽[B�H�yzl~��PP�\:Ei@isZ�Q�#�k#���~��R�S5�`����n�s3�`�#>�<�޾^�<U�F- �^��כ�(��]ŕN�-�e�2�7�2Xy�� ��f�1�A�{z�|	/d�ۉ���:$��ݪ��6�J���{ϰp��H���� ֝���/���*�4��u�`��\�H{#*�j�o�o�����6g�&7_C>�ky��̩pĂR�p:g3�
�I��=��*0x�YS>�F��h��� ��p�Z�O[�;IGo��Sj��s��٨y��P���I>��H�nQk���q�!ګۋk��/�$� q�
T(�C#��K�$�հf���� =�\�P�����Z0 �TA	ʼ�^	�ڹ�w�K��ӣ�����Ä��a���	�������#3*��/��W6b��	h��@�B��C0}����*8��˾�C�1��8��(�����ddENcC/@#鞥�I ��&��JVR	��;� ��:@E�e!�}��S>E���t�8՛Cy�K,s�-���t�$�
�7�(����u��&&ևY���ST@V���kt�"���ɘ�j
m?uP��c�!VL��33��g@�c�6��m��#�w���D]w�zFd�R�6��$98י<�2� Sw�a��\�2�h[l �H�aTg3$�ȥ�d."��;��ۻ�;e$��Ӕ��;�7[�E�X���)��U��fA��E��*�$k��A�D�d;(۵d>&����Q��g�r}�_��Hm�A�Đ/���5��$�� 6�Du#�O�-�:V�M�.�"�U�Q��Ҿ1�A��h�8�a���T9Cэ��\�鬌"Mc`���(�~�t</1*�醧s��
\?�7`��j��#���g?��^�2�#���=�{������?(����Jė�:;l���e���>a]����oC� �v�kZ�A Q������ɖ�����E�o|�5-,������D�$�Ƣ����7�h��!Ļ�^@��>�>��X����=n�m~MVGׁ=m�t@0Vm��5��=,���#�!8��)�{�!��Ȁ ~8�,�E2�H���� %=��ű����+�v� ����q�ԩF��<�бJB���Į2�4�g~Vt)�TD��x}E'k���l>h�/<P��b�Ѻ��׉�8^���
t�yIl�#��m�/�+X��k&(�k��,�<J���[
V�{�	t,T�` ��h!�<�����. ��Y�r/�����Z����]sx�~f��}yov+��m3|��I�P5��G�pe��%[��Ft��^��:�#kS_q��^M��Dk� ؍��<hoE�Q�"��v���Z�I������o�`�����H�S��.0�p����潎g��+�Ύ��6�����쮥j�6WZ5"6�.�=N��i;��v��B���[U~���W�W`�>�m��9Ya�_kML��T�~C����t�,��x�GFԧ�Ґ�v4�䚒�?�Ww�5�׃�p� ٓ����9R;A,>�q�6t��R�\���:�m���Go� `������[��0=μ?�i��򅄙~!���?��I�t_y[SY�|p����e��g齦�9����7���C�x��G~�u�.���Y����w94������9_�_JƭĞ���2m��{�	Ңaw"u���!O{������Y���m�dr���	����-f���j8 ��p��X2_���e�݀B	f�Q��ЉA	[N%am�G�V'��3��w����bm��F��\�ѐ�E�gi��`z4Y4�K���R�S�0�:�;�Н	!8Z5y��s��ų" j�6f���Kc�^+sUg�0H¸A!*�d�	k��d��i�_ ;c�&�0�cס"q>D�;��ɶ1A�;�d��Q�o��}���~�I��&Ӈ������eS�W���w�ӓ�KXK&�j�/��4!�S(0y2����|�f�2�t@��s8���Q�N��*FC �����a��y��#o	U.IO��h��l�o�(N�_�����RM��^�Rˋ�v��Z�1ӵ�Z}�SĤ�T��p����� ��ɖSN+���:������yp�AIN�3sW�o�n6�?��tʊ�ݿm�Q�WkRJ�~Fe�ʌ��NǡGr�8�%��ٚ�.|�NQb��"�2�[;�Y�Cjr
ہc�� H�\��w�Z7�|[������T����rЪ2Ra��'`h&.�	f�-�a��֑�Q��U���D��w@|�As��(�r�A�����~�����dj�di��Ū�^r�!�J��΂̏�	��N��x�|�{��n(�6��n[G�{Ma�L��{9�����8@w���Ի.�(4���;8,e�45���Z�,��k��:����Ѐ��R�ӑ%d���(�3����
���e8s#�xmlBc(��-���\"�a�����U�.},%:32;�J"��[�K���T�,]f�y�������7�3A[%i�L�b�St�WX����մƩX������c�>��o��U��&�-Cy���(�����.`	�>���&lO�gC�¶��^ �ȾC�ݘ̭�]V*�^��b���_�a|��R��G�s&�-��5�5���X��'ń��LTq�|�[-��71�d�L�`5Jɧx7�p{�-v�ƒ�r�O�!t�Ė�asw�{�]�#v�|D�@���0���w`�ޠYL��r��*����3�v^���tعa)D,A�gyɜ��ïD��`���es�]r/?���MB/�3�&��/�^����}OP�R�(��;�@Jb�{�9���%�`X����׽YA����j7���r2i9��F��*��An�y2���j�my�hQ��+��6~�5�qXh��S�i�&T�
���s�D"���C4`�>�V�fBT�C�/;z�\9��+����nG�
;oF��[��x��F� �=kق�ɴ�kgx�M�����)���F�GU
�b�3y���A�s���<C�ݖ"}�'�����[ç"t�j��v�(��8�p�ȩ���|��pC�rg�����K�Ho3I�1���Q�L��ND��E��^�Z������?��_��XT�N����3'i>5�ڰ��ZQ]���m�yl]!E}�z��<�'�/�Wv o*�,�e?_y�I��X��
����"kA��%�L������n�Sx����F������v�͈D��0���p.�����(LR�:�YMG��Y׆�����بR�P�����~�`�Wc�J\W�Ԉ"�����]�/���ܝ�����/��}����̈d-c�l��D~�+_	���(�&��Z��,%y�t��@�P�M��k�o���s�I�$�b|�-rR�O����H�:�1}��nr����׸���P�u
$�L��V*@�l�KC �	}�;�O�g7�?#���?u
~��_��W�yDY�j�1��H)r������ƀ�2���<Zn�����g�&YA��ģ(�>�6N7��j��A��3���n߳DR��#g��o�G�|�<�y� O�P\˚���c׏�.a.�_ia]�V�eΩR�C#ޥ�4&(�e,�)Bp���7H��xp?����/�c�7XD�?^��)DA5��� �cx����w�����dm�Y�F]~�����m��]��Np>��%Iu.��_ӳ�?�j7&%�v��$�ew �g܄��8��6�m�Qp�"��+�T�B �u���[��h�I��I{z�2��BmJ�|��s�&�w��=D"��	f���r]��*?��v�7b���"<��h~0,S<*3���e�[Z
	ۂ�6W;o�'�2�\u;�%^�9�����Hvi(�m���5���v�(W-��6;0�v/ߘ#��|�
�����,`���RG��}sII6n�L���ϽÑ����E�;���O�?�b���5 h�mґ�5���e��E���Ac�0m�U5�
��0���Ng��D���px[Q��s�t6�4Y�gG���4+�%e]���);�o��ӮC��l�ro� � �f���-#��b�@�֞��K�+�jG?���K����xW����H��V@��'{j� �a�b*�y�kA��0*�D2(#D���x�:��rb$_z�%��������A��_J�n\�̑�Vb�Rad\���/�A�� ��`q�vވ��-�r�g����{W��`&6SY�:W��M�WR�Iz�$�{ԻAX���B�D\����摗���	Qn����U)�ɖ��q��=ǫH.���s���Xթ�c�	��XR9����*y���Q��ql��[��;��t�ۨ��a�v�FV�yu�������7tj�5�M��\�w���}�μZ_��,�`���HT�%̆lK�h�33�I �#�>��O�rf�^�j�����aYT�&(r<6�`�5��~��}�m�PmGuQR��h�v�/�3>���VL�b��M+�4�����i27h�j�UC����ZJ�]D�G[��ܫ�[>�F����&c�I?�R[|�����}��e5&�K�\W���.�@�4�7a����\2�x_�^'%�:�f�\��T�b�l�&j��SҀ�.���}D5�v�qڒMb�s.1�]cS�w�R��l��1׷���rW�ȟ�op�ӳ�6� �Uy��0��i�0���$g����!`ۤ �����s����-�VjT��%��P������@��:����v��J��U�Z�d�y7��#Y�AF���Q�4O"�=�IL���z+��Ѿ�ҔUH!G�aNOc)�4a�դ�dB.�!��i��|����V3��!�߫���B�w$oh2[ +��eB5��f'e�$o��ݰ~����M&���f3_�}���k����Jlu��Z���b�L��Ϫ-�W�J� :!�l9�O}3+�/
h}��Jn� P�ޙw>�Ҳ̚Z�����U��mL �eӝ{g$>*- o(0T�U��Rx9��/����6nz��X%�K�K�ls�����TI[;���J��Ia�H���S ��Y.��8�T$O��lr���L�(��q��,��/cIy-�B5x���N��Yy���ݠ�~�#�s蝱-�y�r�KA��y�D��8�_����Ǐ�TTY?����\�*ĊjB�u��^�e��Jg�9�I�Z�E����sh�.���&��aG.���߯3b��'����x��}0���G/�<j ]���g͝o�#pB$����e��s���5T��·"�)_�S���R���[�O���s���@.�@N&��|�-0i��Y⥕��=t�mY����L;��8؅ �o`Џ����g����Vb�$i�����<͒�i~�t#��a��"��S%��_л�+��z��%�ZPݦ��a��rd��A�g�pI�R?��	B�'��q����ӊZ�s֟F�����2�M��;O
a_C5bN�7
�#]�֛b��7���,���g�o�P���-�J�3iɔ��ïw�I]�hT�x/"$��z�,גz1��-�N[�9x��*TN�>(�K�3�$�*>��">	�^}/r��l�I$`ܝY,'��#K�Y��};�c��0KCr�NK�C쥓-Q�5�*�;>U�͋-�VF����H���|���a?�s�Q@٘-�,~x�Q�!(��jPxGj��v�s����>ָ�б��ٳN���ڙ,�҉O�eaQ���V��d�+�)�\�K��	�҆BW?V�q��1j͔�H��v`Y�zx�Z��ـL>�4)R����!�.|@4����/��`2��5%e*��Y2���-��>��/�]4�
��g���^�7*�.d"S@���x$��X�&ꏌ6"�o�u���p�hC�ٌo���?�eU?����O�в}i�L�v��k-MO�����3O��W\��d�@�-	X�Hg�vQ �}}?�q�Q���;o9�|����4�H���(���Erbu��+&'�b�3�۷�������yIfL}�y̝�x>�fĳWL��j�7���],���Jhk�~��S9��<5�hz7��0 �<lp�86�ש��0�#c�lT0�{��4-Z��VG�s8q9��uH��;/��L�����P]B��r�Nm�A�s�9�xl)��.���^�*�T�;	x�ܔ�,E�18�k����65#D��ƨ#��R�rL�1R�.1��b���<�R�;��>4��3�;��1e�����ˑA[c}�f�߄��k�� �I��4�!��U�<d2hi�5��MX'�k�l:����&��!��}�&�8,�ĩ���Ρ�vqd��|��O�r-usJ�������N�F9=�	�{|B��U����r@�	@N�� P�._�4�l:�ȧ�D&��vD�z*�6���q`��T����m�� ��,�׎�F�G:�ͮ��Ѻ#�ＡXy����kd�>����7Exs��>�}n0�$�]~�;��Esqk�;wL� ������nX�B�
�sLG5�}鍥��cb�y����$�naiJ7��9�&0Ȯ<��y�°�+V���Ć'��!�<�H�[��U�����&p[�@^���d�@�j@�e����y���D�ɑ�j����A5�ӕ���j���f1ê@R�E����Q���TW����������6��ؾ��MX!1}�cZ`( �7b�R�� ��'��(�t��	���͵�K;�P!K�=�KS|�&8q�'��r�Z�U	bP #O�6����9E����H2���������A��k�ZI���K@K�q#TgPONUi ��'K@u�C��߁�?"�'T7,1_�Q�֪h��'2��WZW(ָ��]�>�^����@�V��앙��*F���F��L~�RIQ���˞ڀzj`�d���MW�)`�
�~y.ż� N�p��ݳ��Х��(���0(L�e�~�pP�rF��u��hY��vǀ4w��y�����)�ey�a6��e�w�؈~�)����7֐���A�A��'F����}&�5�7����M���ۣ��������Oo�$�Y������F%�y*}L��V�� �>��"Ex9��@���>4S��Nީ�it;#�AMDfд����"h ��I_�U�ߙ��p�j~�s�]��x4�i�Or�&B����Q��4p�ˍ��Ǣ���7������gz�w����I���=C���h��lB2��7��������L'ngq�S�Y��1a���f�PM��"�rh��}��j�zb�*����=	~��E�Q!xM�}���8�G]({��s6q�b��0%�����c+��XcPJ�$VoJQlXh�=��;d2�h}o�a�ePG������Ԝ��ю�J�#��'֗��3�_Ȏ���d*k�9���Hi'y2>&�j���)! 9���2����i�L��t��l�'����G.R�G��s#��gh�|���	Ïˌ�[*����fŹ�Rӽ-���bIZ��BW_d�\蟤e��"��!�Qa%Ԃ��������� �ne��&��<@������t(��@�����}W��nd��x'�����^۱�m�UͬE�E�5�E�]��?K�r�/�W)��Z�YX��&ˈ��(qpƊoh���w 4��g���)J�s�Uc�	����d��3�h[ ��r��k<�����
�{�֑��=�f)���0ۿ�����o>�����q_XR�H�!��#B���!CԞ]S�~����;�J�W��_,	��o�Tׁ�Y��p��
�Z�2�>C�g��#�T@/�Ol#�U9�s�sY����T��nz���)���/�I�,h%�2[V�ɰ��)�m�Z��mѻ��5O�i��5#s�(#��-�4ɍT�fk	��J"��t�5]�Ho��5���&��,8\\q���1\��E���U;�R����Һ?[fr�`�!�uԳ�a���q5�4����%CR�$#�1�㤳���8tD'�E�u����>�x��:�����Z���T�f�N?K����0�?9��;1�B'�f���=��{iڤ�	�`B�l����2��!�������Z5��&\t��A�?T�i�� c�y�"��g4I�Cd���\o��Bqxމ%�Tqy6!�JA�Hĳ����	M�|EuU�g�:�m� �CB��{�+;�%�z1���h�� b�$n�6hhF�xX/��~������Ü�qܹN7����� ���9�l��=%$���`L�E/6b4�o�p<��������c��ݱ��{!%�IޣK_�6C�&Z��o<�.yh�r��i����鄇D�y �*�,S����v�h���E�Pp��/�<��*����l�Ȃ\#��6f+���-e�|�_c/Ɇܫ�q��R ��`�h"��t�jl��?�1����\<3 =(�JYǜmCl�w�I1'K4� ���8{�_���'v��'	q�м;��.����a\�69���|8�V���կ��/1�e��t:ͯ9�u��x~©�,��v�����<��F�?�ۥ��Ƚ� ��Y�Vfz���g���g�E��
�Ϊ	V
��b����cu��qw�T��l�Z�����)�w�!��}U�4��$f��QW��]�Ƅ6��uЯ�I�w��&ẗ́ȯ�PM��w0�km:\jܕ����u�!�[�U�(��+� �6��8r�ӆ}]x��/7e��g�,��,��d=��2^��������)j�A9�~z�$��"�;� x��}ߗ�b�����-���m�V��t�Ԏme^�'��ꔟ�剤{얇��Ӷ+��7����M\ ;�Р�k�V���*�.�;�y������:��/�h��e��iP�ԂtY\��b�׼���P�J��<*0U&�NS�}X.�U@M�{�<��f(EPCvN�?7،��-���x�`z��py!�gcq��Ê2�~�OC��0M�4�pr��k䐊�b���y�ߖZj�wis��fj��U�T��+&�#�^��l�2�%�q�8�6�_'�ʷ�د�ǥ�7�X�V�~)w4�����>�c�)��mzI���:��`�pʋ�jCo�`�ؐ� ���5�\u*�)�2��;}��
ۤ��rp�r��*��.s�r�Y3�L��Ĳ%�"��g�;OIV��z�k�R�Z��䛃w�eZI[����譛���X��c�*�P�1dp´|�j��VY+8�ǝ)���S&:�qE�[�{!Wqt�����ClyH������?Κm���ވ��M ��.��vKP=.�V���k�ii9�w�`���\͒��u��� ������ �M����X|��%�s4賬��C���*�S�i�9���Hp�D�˂�sZ�zX8�f[���^C�F��k�Mܝ���J�ԅ�m�2�_ٞ�'<��tt��ی0�B�.�B�T5f��D�+���X�E�(��CI�8�b���*�C�7)@w?Yh;���N��,��	[d��n��-���S���W��rp6�a������!���oA]X8N��0�9n�7�L���(aT�D�pL�i��G�)�{޲Y�s ��4�L��5�X�����E�� �Cl�j�~>u��N�f��!K��w�x�_�h@w�(~%�n"��@g���7�<\#8��׍�9�����LP��ڃ�^a�H��Y��)o �� ��FC��{F�e�?�9�=��&\x����|�Rd��[�wji�}t�2�S0�@q����O���c P����k�H�s*��<�_&Vrm:Y=`�#�xo/�U����:����#ЁQ�q�����|p+|b�l�O��T�:$�H�a��,�;�c�u�(2�U��sKtOR�T�03N��I�c ~%>]��[E�wi�	%o�Y���i��oJ��Gj��;���c�B5DK؃}�G�}h�ÇD�6�;DS�^�u����V�6}"��x�x�� @�JW\]�;�f����o�
_���j�­��ʚ���¦	!�/��@5��T�V���*1U��i��eʻa#��Q*u�r	�qj��U��F���$`�$R�v�چ�Q>vW���e�X��n�3������1���{���T������4�,�؏��Q�;U
�2Ǩy:��L(\����ċ�O��w���$�����ط-H0VoK�5j�&t� ��$RA���b�x�y�D���F��W皻2���B�Ќq��:��/+>yE��r&��H�Z0����Dk�H�`w� L�	i秊��{��Lሕji������g�.������	1��E�+���Y��2� y�9Un�O~����2�ش�/ǛO?ݹ#P�[�t��#�ӆؗ�E��w�v������C4?��v���6<A�&�ș~��sJ���ygi��)O��S�*~�R�U���L%�נw�|pk�HFZ*������J)Ӷ��LS�Ŭ6�,���d�G��$D��*��^�yI�"�4J��xd�7�~w�F(y`�H�Ǘ7%�ihR�̆� ��+�B���<VK�}W�I��lY���´�|��1΄�$$�g�ݧc�����8\��f��t�!�^�J��
���g@Gz��lǡ�?ٝhL%-<x�iOK)q���*���}6�4����cw�����n���'��)!A���$)��� 
�\�S6}��b�8�L�`��?c��C���0�h���������3��'9���%�4j�Ԫ�Y�㜚���_��o�f���-���m+�%��7�]�w�Xn	ƌ��~]�d-��n���x#$L�+��Lj_�X��e%v��0�+s3�ض`�����C���h3���xC�Qz�AH�l9H��z�Sod�d��3�j����2J���ic|�T>H�S�W�~G2�pE*Y! ��Y<�2[��D����v�^2g)��z�aI��b�R<�h�U������Q� wR���&�:�Q0�K���
�ǩ���x"bIi+����Ec�c�힚�}]�A�	Nh���̩]u���p9"���R�ُ
�6�L��,X�aN�]��K%ᷤ(Rl\G��z��eFõ�t��e�}O�A"c`�M�.&�$l:=�[6�&���X�|&IL���d����$�i�Ef����sP�n�!�|˝U�=V\�������x*s�?�����T�:u��篵_	@וGI����tTVr�`��9�����]��F�aOA4��ME��&tV����t�0�C橼���꼛 ~���{e���c��O��*��te.m�2�!��y��h��N� �{�m�A�A�#"��4W#:��`���"���A5�dP�������8fW�"��[��Gr%#Y6�'�uh��v��N�xIS�R˳f��az>b�&*�'H�r�w�=�Y.����X(x�?�߸<��N~�S�F얍2'�KD*����%5ʾ<;��8L<�֘�{��������bU�;W��e�n�%~W��~wFN�ur��3<�	w(��R�_�z�@�\���<6���觹RP�]�N��(t�"<�xr�=�[�՟b�B,v��ܤ#筪�(�r�'ll��T(��� ��ʼ�<�+p�Q���A����e��','7T1���r�����Yc"������g�ɥE!Awʾ k_�t ��C����wS�I�R�́���`=��M���@�H�`�I�U�wgÈ���m�S�!ƈ �[p2e����sx�����n�Hd<"�Yp�o�myGj� m�xA��	�I�x�R�=�fl�x����Mv�F����WWMeΣ}�}�V�lr�ƞ��2���7L�5�"-��W��)�a$]Os7e6�  �笒�R��'���>�� ƒ.$�S��O��=+V�eA�c0y�3ź��ر|Ip�a:��	��n����)�3�����2��n�4/�o�i%މ���*�m5���'���=#�G`�RɜO�;��E`�xI���AM*ʫ:���fNـ���,�ۺO�ill�i�m���b.�Q�x|WA��>:(��Uk�V��N�����C�\�]��4( Ԃ!䰬��ڲ�Q�z��� �����.�8x�E2qnZ_K?� Ŵ���v��!�P���a��N2s��x�����/�I�~��X@tD��c��aZ�<K�^���Aa����L�� ��xvZ7j�
���̐�����B{䄺�o�&�^�]h���Yu<~0^�:�i)�R�`�_��Fl��a!$ҿ�˵ۚ��,�a�K��u���'��'���[6&-jt5Wn�'Pgxs��2f#�`� `��x��Ò��o�a��-�,������P	JG��C�`nPS�h���]KFU	�>m�PZ�.�ڧ��:D�hZ`̤�~u��|���&e��v�;In{�����?����K+�H���2��Sg�@���Z"|����. �g��(�}��H���5��G�?>�ۿǴ�c��'/m�B�C�����Z��AE?�T�x ��#C�A�=0��U���Av�\<>��+�����CK�v{���S�bƝ��=! ��G��E��J���d��������I�ad����*Ke�u��WE��z��~��ӝ���M�Ɣ}S�r]�����Iv�!�������ꦮ�"���'p��B�C���K� ρ_~!���\�\�E�A#�~!�f�oi�O�(ȐSnǡ�PB��~+����N��Ϭ�d�g���Fe���j~�!�/?۸]+㈖6iA��~/6m.f�X����~r@�N`Ho�	y�m!��5��U-�;�x��ʿƦ�0�[֖��O�A�*�0Ⓥ��w�B�N�ؤ3qL���50<��?mY)~?\[>�?���mZw.\��>Hl�q�
=�buؚ�(�xU=�:��G~�d��	1mM�)I,A����Ɗ��4BSK�IDbs���n�rV$X� �I#�E����hCKMF�+!XB��^�������8A�A����'�J�s(�>N�X��˓��}���d*^x�I���K�p�?g��v��J3�4oֺڋ���Y>#�- q���۱�j>a.]?/� "��+*�i��lVb�s�w�Nճ�d������J��X��6�{��WbiMg6�(���R>M�� �N��Ѷ�Z�� �n�A��E�ZDh�'k�σé���`P�+˿o�)�΅P��\zW̈s���]��v
�Xŀ���M�C�9h�e�1i�W��n1Mql'�#09��ea�o+�χ�}��QO&�ܹ����J��<���<~�/¨`$C~dunWeE�Χ��� 5^�'K��	*����;�u��^�*���N�j�K$�
�P�ej�t���cV�>��oyٴNڙ��$���� ��'�xLZ9=j��*�TH����V`	>�K�:���c�14�h�	mm��J�`\�/5�]X���)[� oO9;s�	��O%��]�������ʀ���;������V$qZ7̳���2���#ܠ��7C8�>#��b�?p���kL�h�c)�@��Q^;��|�<2��î^
GQw�#�̍�ުu9p"�V�K<��(@p�B>� �t�����H)ŰA�o+s�7In��|�˓�9��53�*��[4�ן-��,�����;�1��#a�T\����� q��RI��P��>ӯ<�Wi5��f�>���o�z�����)O֕���
�7�7spD�� ��&�}%���6���LgR�2g&���M�&�	�W(��_y�UH.Uϙ0����+�J��+3�&v�ߍ��S�2�=1�����Ѱ8XZ�v�0��YM�2�#��ߛ���VM�Ǵ�Yo��2>a��[<_��)��6x۷U	���glX��ŵ'�����G���϶(^�+�Є��]O{D$�mJ)�	�Ȓ\.Y�{�ai��7^$1�jj����ض�%��n�!���}H�@�Yq��W�UD$*�$Jx��������F��vY#�oȘ�F��)��a\��-'@F9Eˇ������ V�������`�:�ڝ���ERGɒ�ZxX���#��� ���%�'�z��k�y��&�I�8�S5	O^����?S��XC���(�����56ŝz�2gp������.��+�S��S���8`p��lO�>�0­�2��F�s�fb��s빤=M�_ӈ5#[REٽA{;�{:�Ѱ�e������TS=��r�#��7���n��Mp�a��b���9Y�Mm���w���}�CF6߸J��v��_��ƴ �d����*d�݅Ï$�(���1 ��wa�9�̝^s�K�?by\!����_��M9����D������BUL<S�VF|N{m����R�2� ���$|��L�~�,M��&��r�c�m�o�%XD7!:��0��v���N!��+i�B�t��&���e"Ȁ.s�y�8{�W:t�D��ጟc�&<^v��Ǿ�H@�+c\�4(vv�H �,p����mt�@y�)Xv~��"��y6��]�� �e�q`��}���wgSy��<̘�6�oHP�4�q�1i)����B©��=Ҝ��b����ƋC51�0�=
�� <0��(d@��3�@&�$3ԗL�sy��R�Z]\Ls�ğt��ڲ'yB8�ߵ��Տ+���\w�B��O�!N���܁�WJy/] XٿF��amkj����tP��x�R��dp,f���v2Q�ծSz
�V!�s���ʸ�+2�?=��W8�p$r�Dv�Iΰ��h脒��ԾooB<'?�L�B����:I	��pw� >���C�)��x��}
r�X��`����;k�g�tLЭ���-C�����}�UMι�n$��&w1���mpрXy{��qr�d����	3���/u���d����%�����J����m�z}>���$���m{	��ֆ�{R
��'g��O#b^�n�X[�������,-Sbv~'1qJ(�P�/%����{��]؜m�⭗ޏ�/�-��F��>���zn]�<}X���rG�k7��?jM/js&� #M����H�GKt�gaY\�D��/I�g�}��ۿ!l�106�v,�P�|Q����߅�KA%�~�\�n0
Cխ���J�bM������b0��˺�-Ƹ|:q0��`��7#�0s}4 ^�y)�	�=�S^9gf'q����q�}�����󽓆N�{��Y�p�
�ɹ$ \*����H[������*9�u��wO��tXI<���
��'�Cܴ~�;J���~|�6�Ɋ[Sr�M��>���Љ��E8o8/�-�����ʂ+�H���#,� #d�me M ��Q@)�
(������o��ݏ4�h>h��{J_~r���n�h������Z�*���+�W�뜳G�A;��+����D�Ǻw��Oq7��[q���/h�_ ��`s����z����I�l��%�����OF�ThE6�<,�~��ˢY|�����Na��nS�.Zfk~hʡ�p���4�Tn`��l��Bc[x�]OCQ+�,(̀[Gᐫ����m�Q�w|��Rru�Q6Iƺ χT��!
?�8U*�rݩ �$��c;9m>v�"2��tr�(Z��	ΌG�0U�J����~`;x.�O2�6a7�:[�>�Q�^k�1Ѥ��G]���|w%���┹N�
u-��s����(�Ӎ ���GZm �𥎢
�NT�@���y�8�r�ǉK���qÀ �1;S���&^�JPc5q[�LzFr���x\r�o�O����&���SͿiŦ����/�rqcm�#$B�����a��n:3zʼ6�b�+%��/y��L\7�G�6c�A]{���3)	��� 0��]�y�cè�X!���D�χQZvG�!G7�,TN��S��T������ߍ\����`L��M���m.�î�F9�a��Đ���=�I�s~�9�+lW��u����^�$* �x�"2� �}c.��ǣs�~����Ј*Y���چ<âQd͗�.������h�;ɱ���`8l��~s�Q��m�x�D�fƅȵ�͝ODy���+"�¸�b��bef�T0���,�b��J�ձ)���w��6y��$4��av��qUG���X�P�b0V��Q.�zb:�ː�ƅ�^dB3�Ĺ4!�-f��	��v��o�/Y�l`�ay����Q�i�����$,��r������&oY�2k�HtzvV�:��@v	��s��{�ѭJ��&t;%`��0�e�*���F��创�[���w:>����	,X���L'�&~κz/�|��'�K�H�Z0~J�)��9Ic���-�9lI���oˑ��|��'�h񿩆�s�G�;Lu�	� Bp�/��Ĭ���R�6��iڍ|��.R�ͨp��-2�S���a[�����z:%"(6��7����M�SLU¡ړ�N���0���K.u�m��9�A/�R=J�4�T˖H��1����4�#�L����{_��Ur��Z��6�JFY2��2�%�
&nM�]�Q����BG�����Ÿ����v௣������9nv��k������[����(���6��������6�?Ů���~/�\�βۄ�
J���rW"7�F@F:�*���/�x�nPmФ�$ls��6q6�t���f�����pXi7*����nI�6_��"�xz�jYқ[�C4wb��e|0�G"�+rQء����j.��YCD��mח(�R���V�ӳs��o�IR��jޚ�TF�բ�*fg�=����#u]H� *���P�߆�a��ЈȔJ�����>�V�Õ"�ogm���P��zܥ	��X��+����1y�A	 F�NG��9u�����]��KG|v���_�T���Ѡ߽�]��C�̃?��:'U��kP�U)r���ǻXH6&n$��hw{���(*�j�s�\�Rxi��lYQ7Q!fBr��L���3W�*��0QݜS\8$�L-���|x����{�*"��h����x;�t.�n���D�?;��49���t���w�y_r�#r0ByX�������@�_�&+�I��b#Z�:�$t9�Ą$��Ӝ����EP�"j���9>��{��O����HKS�&*<�	��R4.����ځ�8�����T��$�"'W�@1ʣ(�$�}X5R��Z�.�+��J��ύ��0]0��<O�c�^M�o��S���D��7ǤR��n�_�1����f�F#�-�4�9�d��"i7���峣#�Ȝ��(��d���:��
?����3Lx�՞���D�����#^����)S[!4�Q��1{��]���ޯ�f��>�"��V=|��1�Z����p+�UE�Zn�S�����Yb��b�L�1Ȓ4zR��plϋΈ�>����/s>���R�����_5���>��8���j��*��2�FD_�J��N:.�,3��Dcp�g��s��9
�ҽP5n���[��"WaF��bń�����!(un���FR��쯯���a��z�AJ��r�^�G�(����?���0���O��L&>��_�������0ɲ!񖄟8D��@��	�Z�wC�wð�q�����ٯأ��jB%6��Nb��KMA�L�-@��ڄ�D�赊U(�6�&Y"o0�uB�x������`O6f��5=2s����]���0�g1zn�-�(�e'������ 7�JYR��� �x���h���'qF��v���d��n��1:0XMQ��_W��T��¨k�e~�{N��i�Qg��F�;��
�FJ��[�b�ՂS�!H`�����P��n�?m�
�
1�܇��hMA6��#�8����N0x� �G>Đӡ �#|�� hD
~�Mgؼ�b��W0=�/<�-%$�RG+�1���!�(�z]B	�{.�_4��R�+��D�$)���D���~�*���R@QV�͙� VKÅ?i��c@ N�J8x��"�Р�IW�Q�������"��wΦ��d�d/�)�hI{�&Gn �H�J���׼g*&G�T��w���٨�.d/��5��u5��P�$��>ࠦi���8�\D��s7��c!g�W�"�x~�s��������t|�f9��xU,s W�_y}+Ho� ��Nsܲ�F
Yb�6��k���eԋ0N>���W�sQ.�+D(Ȫ�	�a�M��y^�.N��"��~���,1������Ѕ���_j�?_GR�fX���� DJ6�JC�}U��E*X��ϥ�=������P���?���� ��Z����F���?��&0���<�%Z�V�/������Xl ��UCp�,E�
5�A�N'w�w2�Q���E�6R��~�x����W�L�2���D�R+[J90R��y�
'fW��gj�Imdf狗5sYI�	�x��lu��\aUJ���U���F���-=��*�S���*���o|�ʆH�1p�Y�����Xdr0�Rj����x�yMٳA.����s��f����,��fԛ.���=m���3�[%��xW�(�ɤd��ψd2T����A*\��
��s�q� �ѓ���_l����3�*��q�E�_:pFF,���/��Ҋj
A���w�3H]C����𮁖S����ϣ��	���{����ɾ}gJ1;����9)��L ڃ,������W���~����V�r�*���x����7�n�Ne�jH-�M`����:��
򽨺��Z��g֊�yMV"��(��f��=n>��w��!�<3�Η�tԘ��G����_~�T�AA#Z-ǯ���(s[�T��.�kz���n�*��]a��i��h��ei|�kz�;�a����O�Xɢv@bT���D� m�t2TXλ��:����8�Qp�r�����A�tَ�hI f�M �� ��IE�8b����u��������e���`f���3��^��?FD����]}:��O_���:�ң�m���h�*�)�Zz�������r
� ��f�QC��-���4B�/���l6�ܒ���*+���7'MZj$�.���R�ַ��nC��f�rk�ɜE2���$��C@E���l��<f�q#���M�ޮ"ڡ�2��t"rN�B9.\�g�a��k��5ht�x�W;PӉ�h�?X��B�곏�JZ4\ �GO?�Җ������Ҁ<2�����N ��	�t�t����B]Y;�E��g�����Ĥ��j1է�f��eb��̾��{��	�S��_H9}�]
� X��E����@��Epa��[�{��?}B�@����K��c�f�r�k8��%�܌�q�q_���Z�-�����V����{��p�̓��2"Zw�:�(�i�/F4Df�
�2J�m&]����#�64ї��,i@��G7�>�,��*���N�:�ٔ���8Jg�xP5�d2�V��gQf����B�K[S�J�u�s��v���a����vt����i��04C&WJ�	�}������!�>'�Q��m%%�>�� ʒN��YC��9x�Vp`@>޼���j��-ٮ��X�T@6��XxYƨOo���G�ӹ�qҀ�?	���5L؊'���#�}(��|[��:V�@�l��a�*A<�����.h	<C��y�;��6S"?	��:��sC����RQ�8K�k�ĵF�?�^f@Qy�|,�`�S�����{�t�r�����z ̟2��R��00���1?��*�6&	yƋ��=Y�c��!g���QS��)������5k�Ƞ�W,"c�Gmj���\�utP�/!�]o �A0�燸V�w	u��b�A�4��7�H�� t\͈7Eφ�pyF��c߹pc=������2�9ɗ�]���@��o����9�!����p�n����8=M����SiD��R|kv�`��>s��͋��
�z6��
ەQ�N��k��������l��x��VE�9��l��8dCmʅ?����=�^����m���؃
��?��y_�`�}���<�RPM��$��
F�
��E�����yV�huq�������>  ��+����n1\'6h��g`G*�t�����=.�6w� ���vV�/�p��aS�(��V-�=�MA���8���2�q.@*����I(�P�ō���6(q��k���JD�~N�*��o���*�@揽DӖQvt�R��Q����p6=
]�� yܨ��T"�G���'�y;�����2\� ?:��<m����h�i�`��rF�����U�0M�r�ʁ���[,��xk ��5��m$��g��L�GvN�����YWf��H'"
�����f�I?��T�/�Ԥ��zߴ����|y�x!UV��[��̮p�Ưv���a�w2V���OU(xg���HO^D(�Im�ot`j�{�����p	�����(��kE�(��u����D^��g�Z}�|rwϢ�)eQYw��@Z7u��w�P1v�u�ԣy��`��$R4W� [JۿD<e5m�n�CG�S� E��Z�o�<��V�QLk8d{��a���o�m(f����:�����t��9��C�Cjc�h����\� ��/ܽcl#�����i�AW��~�B�Z����Tf�}j#�Vk�b���m%�sy W�(��GM����ҕ�1S_��Z��A|!�Z 6$���$6Q��3}^���r}��xA|rD�,�𷯑o�^�2�T�h�����"cC/s-�(��lIկ��{�̨���-x����A#��598�����fU��a�F���]R�#��l��ifx����eF3�	�u�n_U&e���'5Ab���q+��ᩃ��ՙa��K<��0�:6�D)N�@@��ӡі$k&SS�7B+��|��](�2eҘy�'L��,�Fqf�<�3c9����礤�,k�6�=��(Z��U�KY�.��89w���m����mr����f|��Z@����s츜qȧ�p�o�S��뇂�kH���3_)b�Ku�U��z^r=��?u���c.=R�Pi�]�$�x��Ć�&5tk�[�ÿ���m;�Ր�B��{�w~�Km��A�(iL��Y�?D�V�xyJ�m�f��>��I��幔|���/��1z��p��4��[˥(��^pe���UW&fa	h��Հ�y�V"�B��8��3R�]I4�M[M�De�۫�1 M@�ž�5�}��ɟ��\<iܮc%��*Cw*�`��Ѕ�~��+[�1ox���,����m���pB��9ZX���*�ؼS*�$|���z�8ZR?�HO�f���J�`��4���^�6܋�l�C�#�.�Y?'�Ú��j�P��B6KEr�۴}���V�悗��>	�5�� d�b+�Zu9v1%��-y������k^|�ޥBy�\�U�S ��0ס2,Ƣҁ[�	��"�՟f���d-�F���_y���C�fq-�M�n&��>���	E?� |$>�xH"bcr�XɴX0
#�&�-ւ����Z1��t�,1�٬�s+|�+�ո��0�p��%�x�	,���cC����&PiJ�Q]��6�+�P|�SÃ
�I�k�u���,�0Vn��]p��L���V@|�^5����\樜��(L8���Lf+/>p6^�w�����9o��c���K��}ig��Q�! #{�V[*z4�����W��N�
E��<|D����&;��F�����.�J�|p"ײ S����>��l���x:�4��t:uư�!��7�+������c�=Gz�����q�̛�$<�A�_�E�.�P�|���鲼_B����t��%�����x��z�:ϫ�?^&�	�c��|�|߁�~�W:�5_i�U��!,7�Oe�+���`=����mЭ)�m��m��_�R�;�D�{]-�@�/�rd�������=y�o000w� a�,���p���F/��:�ɒ1����3�[����4��:�19�D��vP�>�7'7�Ca������H��_��f���{˧m1g��uf{��p��ZKiG0̿�V/�
�s��G6�5��O�O4v�,����:pR�K/�`�$-����Y�����q� Kv6��2��������B���J=� 1AR��a	x�I�phB�{
"S��Kk�Ӊ�K�R������*��^�FXn�J����)�H�q���֑KS�����Nv��'��H����s�$��纗�7E����}�i����:�vf��md҈��K��J��s*�?� �D&�G��d�qy��R<)C2��.C^?�ӫ�QtEl��P���8��;��Oռ��>Rͼ�6�q�vL�i����6�������B�hP훾�,/�Q�G0`u�y~&��"�(�q�	Sv�)/y�K���u�y�*�g98X�j���j�[�76DbV��t���W}٣yob�m�ҧ�+)P�����q�z*�Y�"���6���$��jM���%���I�$��з�*����m�=4���@��1��	CEC�M�
@<���4�nu���������sv�}"X���X���,�	�/�"��ْ��cr��j�}R�ӿ�k�"X\O�1�q/t��{c�������_������	����9�~׋$+5��":J/ʨ4P)��VA5��kI��[�3E�gdTx��D�#�Vw�X�͒a�B���ē
G��d��/�+�rl��~�aM�Oq��0���`�ݱF�J<v��u^���܉x�C�Y���q��Rs�@6�E��Z��w�`,&2�B@&�s�������չ�����>�V�=Xx�SuX?��I���Zz�t��4�奤��Yj;2���c���L���"��9p�o�������l���겣W���A.��eD3:9�}��D8���>:[��uR�TUɥ�L"��.��b�gQ���L����l�۠;8�Vn�=�ɉ�p��cU)� �h���_�;�~[X��Ja�/(�?�V�N׶¦X� I�MD~�hk�ᬮPa�H)��������?��j�=`���%(NH��}���w�e�;K�7n�j幠o��(��_V�r�8�jKOi�En�ȹ��&^�b!_�U鶓#��i�l�>Ԇ�X���ڦp+Ϡ�+W-�ڕ��_kU2���N��*O�6�5R�s_j���Q��WI��0�<*ĝ��3+�8��f�<���U5�BBk��@��zdx��*--����1D0,k��s/ޓ9#�|��Ro� ��o�a���c��ţMXEx�F__8�R�|��5R{��1��]�⓼� j5��Wj��������NI&��0{7�F�8�#�2�$-���$['稯��+�_�b.(�=�(��K�$��3�� f���G<OZ�^[c;��nMq��CSj��B�L�^�4ԡr�FBp_r=D�vHr:��.@��F��p'!��P����\�-}����^�g�KTYU
���S`��ŗ��g�������-!C���B4UV5$��j���(y2�ٝ`Җ��3�"�KH�v�8��~������K-_$�9_&�u4�k�W�� �.՜~�R�j����P������0X�*�����rΙ �<�ʹ0�WG�?���'8#��s�G<�t�إB�m5��]I_�v�	oQcҕ�<1�!6o��ۆA~Cu�:��V$GUJ��z��/D6�5�zr��R	��.6������2��&�!���9�${��D���n�!�Z&�V��yD�g �l{���{>�F2�d�J���I�=��d"3M��|*|��
QZ2�n��5G2w=E�"�Z.g�o��=([���D���ry��nQ4Wۨ'o��]vCPF�lf-�w3��Ig5
�c���!ĉ�u��u噾�C��[���e��K"�9����O����RWV ��m%�/�'�c��nxJ����Rʋ�9��c��7�5�BfWp20���E����2��j��M,�!IGX˼X���3W�(�|�=�q
OZ����:����E��%����V�#ђ��v�C	��î`�h=����:���ϖ���Qm1ֿ��$��S��M{9�V��e>-���ϕ�h)�pX��mƩ��N���Id�`�:��+X 1E��̷�����6����PR��6j��~hebr��vh�����I�r��� .����a >�	�xڟC��m7b��Wx%�\�Zʻ(�i+��4�!�#o7�w�nG��`,xW�����>����9_
)�G�g9m,�U�
�vY���ˌ1S�x��:�FL�:_����$���n��" mN5c�H yN�S��#F~Ȇ����ybk'^\1�=|T������Q�Bf��V�HjȜ{%Ϊg�k^Se@9��D����@��[��<�E�:�Ƌ�:v��]<-6��'��(t��>2��S�:�^��"_ȉ��@�mP�y�����|nZ+N��ei��"��o����M���M�(�w:�z���,�1_Ř�X`�ڻ����C�r��"�`� �yc/*=��z�����v�U��oS�q;b����9�Q��A}v'E�_�1��)���iY-o|T��;S+���P�~x^�L�3N3e�@�g�O����������@�A�1����.�"T�v�;CD��{MF!ԧ����0&���cm���f�8a����N�f�Z�jӆ��֯@����b���I$�T(��T�tI��i:_�픠�X�o�d��#FF�iɹ4�@[�!zN��=��Γ��n���{l��+vm�$(�a"%��hk7tKa��� 짡�ԎZ/n���r������C,�a��c���fR�T��0��z_c�����e�	���``u�Vl�9�!���O����ax�2]�X(���o$�_wnk�cZ2�5v�AS���*���,���{Q�i�%�� 
>�K����( #F�[cFT��i�C��dE�O���'������T�N�� �\��4���K=kc�nv�\�ړW��4�y|[�O����ʸ�
b���!����e��.�10z�X����'a�]b�I�Ug��t�1��a�r�0.�EGך��K���	����>�Y�h��h��(�.�� �C��� X��"P.���XTOo��}ͽPK�����5���%�;P75�-{*.T�j�����`|�p۩��O��M5�Le��[���W���|��ոl,O����%//��| g��:vhטV	�W��︘����W5~`q�����Ov �����oHP�m�c܁)�_�������0H�ָq1��|��px�b������N����J��~&W��i�g��U���r�]�fq�|[��n�0Up��`��`��Rf"՛���جm���;�@X]T%�$�4�h)���x⾬@��{D�u��vD͆�/r$tVf����R���?d�p����߹|t-��4���E��z}�����>��a<*D,$�P#[o6~C�T�8��z\�r�ڂ$e�Fd{�q��	���3׸�����CC ��!eD�&R!��OY}�P��{`t������t ��a�X��H\F|�)럋�7*�Yx�U���!0�(f�mx&�m|i|mo�U�볒�bP�-������=�k`�E����9�2�����p)����#� W�f�0'�)T�Β1�$��pc�i`Z"-y�?�J�P��]V��	3ۄ�Z%q�����Z�ܓ�cb�9GR$Ҥx�/]z�DyO����ӡqix,�-��R����w�|YMի����(�pɋo�YSߦ(S�֜
��d���k�OM,�w���W;E����BC���Ύ"�:�|`{v�fb�@V# �N����VzPrZ��R��u�W��tK%���W�\�D������$|2��@4F_�-=�OZ���z�ٕw����W�+�Pk���'�w�m#��%�Ɗ�Z�O�\X�V(���g��H!�V�C�.v������O��gÞ�)m��Auj�=O�r��}T' kO|{�����"M=�p�;+�l�ښ��,W���Xs��'��]����.^&@_�}� ��!v�;���܈&Px��'�C�A��Sv�:!Y�j��53��L��#��JC�p0�M���A�]N�v�����6	l��	V+�cbT��S&v�ADي��#�Ww��<p:�������m�M�́RM����p�������DP������A��h�xm������h:�>��ܕ���ط������-�?�|���d=�S���n�rx�Ψ$�#m�-�p?6��� �9�	O
D��x�@���&f������`vVFq�m1��	����5���at�?v�Lr����ʎ����5���i[����M���	ʃ,��N)�6�U�a���UO홃�f;ʹ�����P�*���}�,�{x�C�{ަkػ��k�`��P�9�i:���,�o�����eR�>�a������1.��(�}Xm��ä>�{��0���⛙�{�Ж!fV ��`z��4
���梋�)/��]C5Yz;�;ÛY��������ur��[o6�[I�ž���D6H��â��kv�)�	�$��W���QlI
�P�~��l�c,�犭�΅Hmj�,d(��4c��*n|j�ˢ��XT�v���4Q��w�F%l���1�8H0�q�}�^�)�|�p;���T�R8pϱ��B�N��x�e�Ǿ��w�l�8���
��4Umc��>%`m���;QkMgK�r�#�����'VJ�HB3�R���8��'᜛T�������~f?
&ʵ]U�t�=g��f%h���K蛱��_�"��,x+C�������g�pNL����V���[Ѻ�\v�����=���K�ES��-�,Qb1#�-j�C�8Pv-�-�U���(���%��ݤ�
�����a� #�U��faE�#��ҝ���K�Bni!�E
��%�����u��wG��� 8c�������3�X]�x�8g�dGːs�[WN�J�,QlOG��#��t6���[��/�<�dl0Y=���3�O�y8��a���X�L�h��]�ʤ��F���?Ѭ.ē{���8s�▅����_]���ѻ�J�jl�����^'�zKc��o��N��pD͠8�\�f�!��X��I�OV�N��o�>���ؤ�\�l�&~C/�j�d�X��!n;]p���/
�ؚWF�b�ד�#�����"������RM_���[y\F�IUC�F��SK)E��(A���᪼�s�f���`�����5;���Y@��_����e�C�64��!Fv,����Rf����"��L!g�2I��4��I���h ��#�Z��,R0�~�1&:�j�c�GU���Pa"�Qwv��}�9�N��_Y�+����޲���W>��8#r�7�m�Ԩ;��������2G�?ύ;����[P�tޗ<��~�g���Z�Y�F������{}Nt��Ӏ_����_tRy�*�ٯ�,�GH>�-4$�-O%Fd�*�2� ޳�]��x���H�h�����Ԕp�5��!9e!,W���j�I�跋���QgQ���**� �;e�,�����\ٔ�Y$����=�0*Uo�ɮaaO]�DLxD}L����ҌG'����3�h�P�W�ڞ�X��m|�f,�s&��@��1�`mؒ9��J��Ǳ�~%�UĖ��$?���]�c�6Ll�nq����S�9�T�X�<��y.�~�V�y%riĩ�&�*#��nq�:��"������ڈ��ciA=v�Z*��|#*��2'6x��i�\���ȶ�+���tf<Y���{ȋ1�㴑�L���J�L��)b���,�xb/M�+�7C�|�����=�V���{�A��W�Q����D�� �{3���.V��#C%,ޯ���s:��K��z5���h�V!ٓ%Ϭ��*����;`��n�e�Wf�.s)��%` ���3�4��;���O�$n'(}U/7ʶ���&�@����E8������[��41���4d<��o����}���I���V�H@�=�]>�%	]�~Yg)��h !Ӓ� �ռ/��_�E��rJ����km��5�R��R��s��&�d�U��?���u�p��A�T!<#ح��ӛz;���.Y��@��r��{���GtȑL��W:3������:�}�׏|�wk-�`|��h>1IV��+���r��uOCT�r����	���-ϖ���� A�S�K6Վ� �����fba]M��5���>MY���qm>��3+
H<�_�������-��u.U\��j0�%�[]Қ���$8hJ80Ԗ�ͰՊ=C�M!ؕԫ�{$�>���s��\�e����Ã]dȈ�^�"h�v�4��B%4ޭ�L���X>:}%�4��WM�����ɩ�_{e�V��Ut�hM�64N��[���p�êw_��ΐ�G�"�4�Wk�+�������Z+7�Dý
D]E��e"je4��7{�J�bCr˘���`i�c>|�Z)�v�$p%x2?=7��\� J`MUsZl�tU�s�j�S����F{��c�|�����X9�m�˿n���^h+\��|KB��n���h��=�g� ?1��E������ᲀHȨ�8	�^'���&,�@.��k�Xz�����2@P"�j��HA}�f���?x�1_%��w-��I���i��ƀ�e����Q�Ù o6筒=��:�N�usy�*�4F�p���cʝƓ3�٠��e�v
)(h��{��87;Gp	�c���;EE�^�xX�q$;���dC[-�h�:�L�<�ރ���+�]�:x5��%�B�:�`��F�rc�,z�b6���`#R�� ��yU@�L�j?�p5�ҨU������L������X����I�BY����z�F�B����%~=,�C�1�e9�%�I�T��MM��`1f��\���%�����9�I�� �V[�ٌ�zC7ؿ�&�<Ԁ��d�dQ+�dS�͋���R�	"��a\�v�ǝ{��M,�$f���=7�8��V �Z����/.=ɯ�L	K��W-��ڱ��HL@z�[�D�)�q�'S�_��T8Y�/�wӭK�	h6ubB��P���T{	K䤅l4���&<ݽ�[�H��G�ҳ/�ki���خ7L�I�URr��aus�7��V$܇!\k&+�6��ࠟ�J#����9�=*^�CPJ��N�ݾ;�d���u��F�8T[�{�Fz=�w?��P��wH���e���%��x�N�>�g'�͙_s}a)�CN�.(Z�t�9�����D8Mt��_R�^�={@�@�&��2\̢N2Z�&d/V&�����;���8a��#�
�IX�".FGA�<똦��DY@���|�(���'ĺT����2֨�l�1�tS-������0ګ�yq�/?��MIh����e��5����6����l�>�Mc ���6ꗅ��׽c�0���7���V.�A�NN��ۼ��-�
e��\T�@����)�����g�,Z���f}�e�I�~���&�V6��Γ&�`�O�}7�
��;L�q�UЀ����&(fz�5e�����_p	�ZQ�3���y3�Z��ea%0/�a��h�~RL=ƚE51v� |����}̨%[��.���Wn��<g��P=l��3j^`���NX����`���.�e̓�J�JR���}%u��ź�W�	0� ނ$Yo�>V�5)^y���qg��&k7K��!�>��J!��">���:� #����=s�hsO`o���pI�n<�\�d�3�����;@Xl�Ԥ�_[��(����K
��S,�J<g-�.�Al`(�����d)�c_B�
��y�@���\��ގ�}�z�דt�PaW�w�_ܽ��e�_�=]_-A�e�_�U�v���}E��%WmTr{a�9����Zc�y\��ܢ������G��O����A�^ɘT�O[kb��V<�&�$̌^�`%�� )�=�{8
(��M�k��3m�������r"���w�,�A�|�p%�v�?>5�&��F�*PV�S�8W2뷊���R�T���f�t|�<t�F���Jɑ�k�>Xz?1�N�v���>!m��?�=���N�����d��R�bH9��M'�:�j�c������ƴ��ct^\��'�+�>u,y�V,r��'�<����j������ ȉ�y3MG	���e��Ofg����O4yz�_!J7n��ꈮ�~�z5����.a*�S���i��(�b��ҒT�(�6^�g?��$��!NǞ���� �k�e����� ? ��B.CS��Ro(A(C��-���[c/@��ܐ^s0�GVc@bM��3����;v�$Z=k��T�G{���V}�"?�����h����oy���7�Ϲ�W��:��s��i���T�"#�v���A�J�'!���'߼���������bQ=v��`�����1P�^�^F������C�����D�sF3(��j��Y�O`�$�J��N����Oi�@Jԧ�R�~� >�@�!��Y�&�6�=��=5tS	�pI��:�X��C"��b�M�^D�w>��b	�%�B��^yzYDDH��!ɡY?75�����*���ạtrÅ&� ;��X�!��XlW���$�c8O��d�@3@d)�9�T�Qw.M3�S��x��k�b����ZgT9Sa\5w*�J3�'Ӱ���Uj(LV�e:�	��>��<р#���	L�t���Mګ�����M*ƶu��v��`ۛ"��W�*�`�(� f����9g63ǂ�f`��q8�yYq�|�ఈ�.Gaygv���}+iŔ�RF�Y�eC��D�Y�z���i���fy��"���n�O����K�_�V��d�9t�$���o�{4j��+�@F O�NBͳ���__f�����6='ʓ�Qo�tˈQ�t8�-џa��3�@�ߥ;^f�R!���*�^ܡ�J�1��(7��&bD'Y�Fv���|�l2c���h�����&(W���Q��.��>�x[a����6=��Ӿ�x���G8�B��S��L��x�"v:��c��Y|��b��Y��
ɎA�fyt�ff��{���%B� �3�2�^��g�lY����H�C]���g C9{?������d��]0* �
�o���=��\~EK��J�
���ID���9��hX`�l'|���n���6T3�V?�%[x�����ڎj�_� Cy�E4��C��h����<����眭��䶣(��6�̱�K����LmQ��l�te#ox�0J��33qn�� ���f3�h�����vҜ�V��	q��XM1�K�lⶃ
&��R�F=��6[����b�0��UX'�#����?��;aH��}.�66�*����L��[����-�'^���k�8���1��x5��y?�WbC"�����*����N�!ɶv'p�Os�N|��LQ1��yZ�I�����=>7�$BEkn؏����-�]�s*��ᵆGI�{g�|���-O��]I�ZO؈'5�g�n�|;�4�恮�rxh�1ݓv�b��(.o>'HzV�S芾s�.D	Z1�NC���~��_.r" �GP��z$a�Uխ(��|�Q5L��������y9���44��PgSyL�(&T^�)8�k����#-��tbz�
���ɲ��?��SND�#�Ėɰ1�<�Mׇ�_P���m=֪_�n���̂1���w��� E2�G��N��J���H��r���
z���vn�5�0Ro���"�D��Lzm�T�B`�܂Cxz�p���i���ڨP5ld2Y�Ӿ�&�� c�͞�(��z�A)�@~��r���aΏŹR��f�.M�d�w��E���Fy;㪌�ѵ�R� �m�)���q�@�q-N�f���ںC<^�l�����9�˖�F�qp�3��S}C�.���;s��SYxQ�4}Zp�
�mx�2�M��T�38W�ۧYٸg����z����$Ǳs��~LcmJ�VҐa�[;g�;6�SyW�q4��L�d�N��50�̬�nW���s���P|b[6�!��HLk��\t�KR�6Y��Eᥴ�t�E��:{��]�I� �,)uٴ�z|A���	�Vu�"�XZ�cA�����F�JWg}/p#�k�B/���1���1�8[��(�}�
Q�fM���)�'�˽�t�4NH�)
�.!�Z�E�O�Ӄ��̔�m����4 >���
�X�"/w�Y�6I�b�:pa�6̝������O�<<\�~N�W�� �5�������5�`ŭ������CJxm�C�L[���[�T喸l?e�����W�S�j4#����,ٕ]�Tq�3pV9v�$T��?�=x:ƫ�����[+Oo*�=$�RM��O���e��������'w+�¸��)���&]��8���e�Y�K��6�ǅI\�]�DR��������z���=��[�����5�%�	Yt9M\���ʍ^�;V��P�	�WVL�|�GS����*�+1b�_��b`u����lb�[���1Lܐ`[��[x��~N"�^���Έ�m��@�;��)prwg��I��||���Ћ���\�a.��
i�e��Ó�dl�� ��+r釠q��y��*e6�2P=w�c�}��z����w*��rE��?�(�b}�2�:L��sp��U�Kj�P#'��đ��fj�@1`77��������D��pY����ވ�i!O��NTC}�s3�}cQH=�hb�_	�	T�$�"_���U�B���Py���BӪ��[�:�zR�������:�t�$��8�����>�}5���=��+�AmK�3��|���
��vG_���Q�����_�Hb��~��.O|(�ds��0�T�3�f]�����T��	�R������%������ߘ������+��|��^�o��	/f[�H1`0\�Y$�q�G������ŵ�:���@<.A	%o:ۨqķȅQ�]윒p�����n�f[E|��7��2��c�Mpq�ӱP�YP(#�e���
�ڷ7�s��Z�7,O_W�N>�������h���՞����8d&�z��)\��>��
��`ڈ�T��_�@�^ZO����=bQ�V �e �;"]��9g8���� �+��o� �Pǉ8�����]�N+$����A�mM�9�l�X�:������*�E���-p�,�y���z��U3��E���iP ^H�P�ĩ�o��5���+̏�u�����`,������u���n�M�	��TR��7�f�q����u�8��y��\�����u_�I&�O M;�>�+
�Z�b����6x����cK����O&�7�@����5����T C �^$~b5ݝ�
��rl�%h{�t�hq�	=A�w�k�qN<��J]�?���L�����/>���)���Jw���������I����3J���1�����������(ڤT�B'Z*����^	�*��c����=��dc�^w�'ꅷK�����u�p͞BΜ�;}$�E�
$�5���Vǡt�9�S�I���$2)�m��9������i>x�����>��x>�^�.�#����}��kh^��v*��E3�Mՙ5W`� 1|��tB�zԋCZU��/�`x�N�R�o�3&8=��� �����#�7᭛����y��!��1�O��?�B�@v�R�&g�
H��e��$��qm�K����,�-�W�Oҏ����+�c�Z=�0q��캣�&Ev �ò��ə��dCB���e�50w�Y�K��b��L%<�&C�Cm�������S�h8R�aFP����7|Z�&�h��@Ԉ5▐ι�v�̈́��6�9������|�������iw0F=�?�̓��|��c�ɜ��r�����w]��;����]dE�h������\��|�2�'3��/�i�m��p�R���t���=�S��$r
ۺ�[i��h*��ou���E�Ъ��&^
�e�1r��M��N��@��%d�|�	NGU��9��h�+ˬY�kb��H>�����*I�	�;�s�b~Y����cfPpC��Ԫ^�;|�!A� �+߫R2�ֱ��׵���n�9��P	������/{�w���AUM�*�_�w�Sׯ_I[qL\Pc#N|��9%\q��{.b���k>�$�vXEh_!�f$��>�����P^Fī��ֻ��F�{Y�=�@�n!#]��J(���>�v;����	�>��=��0g��+�Ҡ��;Q��
C (������VJEce�5�����	�W{<L��{A�1�9Yx��LM\VK,@\�aA�=yh�l����H�o����3��Դ��ۖ6}�s��&��;���G�&���r�k����c
I(D@/.�'䚌J�{�9{�*(Y;�lK�H����&�}|��:���@��� q�!��$B2�b������Y�z��ѿ��:���>�nԮ�������y���0�A7߻�f��
���h�!?��N����H�U�<s�|0���;'��<��7E�p�}7*ĥ�����{=&��������Z�|��/�e��İ������@ܾ�2Pb_�]4"���Ԗ���ϥJ����^�$QԻ:QR�?��1�F`Щ�/1��uĥ}ͳ���Y��'c���E�T��D�Pa�q8���'���Kf�>���M��7��4@�ӖŅ*0�G�1��4�,L�4��MI
x)���约GR;c�%"����M
	�����o��8Xa��g��jz�K���5�*3��n�f���%�)E�S�c��R��n�,H;gih%���VBN}�\�A�(K��v��k�NE�w�+����K��������Fi�K���B���Z��K��hQEy�{�$��q:�����*���^,'=]L+0����P ��>��.ݗ3y�_�$JZ�+���E����=��5M���xn?�8n�ti3XV��O�\d
#>�oC�PZFy64}�Cj���?��~��AE��
TZ�̤@���0N��kX�g����P���ՊlMK�G�8�ee�gQC����d��l�.�H'�l�Lh�Tw����G�PUbLФR�2��� �j�q?tR�^�h��غ��ŧ�%��"l�.~:�몘���� �f�>����E��]a5m�u�jN�[5
IB��?}r�X�����r�M|��B�5ړj���г5_j�����^\`�MQ����������m���r��D��0�%�FP�~�K��a[ʌ�z��#[PN�v��U ���kX��������8b������-W�3����Yqjv�1�C�7����[v!w�2��E�/E��D�̓� �X�j4���-D�N����EW!�=O+����Ӽy������E�k�Y����#�+0�����k�n�8w�\k�R%_'m���^�i����>���]��M�ve7y`��o��KDV���b�du>t��TOΏg{ēK��*����O�.�G�]k*
��[J�t��x1;y�1����	�'�;���^PW�!�P`V�V��7���-d"L]�t{<���7>����L^i�9%��g�\`��@���Ș6�T"�Fc����ǯ�mp+�i���P=�ܠիC߻:�g�`�FzPf؃�m�.N�_ZT����|����Ӏ�~�G�-���?/�y-��_$��q�/�s|X�4����������w�vUq^t8[�9�ɔ	��T���]zdv��SN&s ���n�9	�����V�K�Lh�R��,ڊ�s�d̤�ۦ�!ʪUʑ݋1��9H�C���M����~kO�ۈA�wg�1L�+,d����q���j^� 52c!��J�a�f]M�jbD{����u2^D�ɪM�U�,�WU�O䓺{�:u�7L�܏��"<Fz	Q4���@'kCK���)��x�o��̐[���8����#����Eԛyu`�L��پ��}�X���c/���B�οv]`F�&�]{����H-�Eg�|Ͱ"�����W�z�7�#��0�0cSW|}�U�QWX<�KrK�#�c��G	p��l�PJ��;�I<� #G�B8I�G�#4�W@SHÁv;<Ρ�x#�ܚhm\s�W���(.�e��~��?ɪu�%=/���%���s����c�������6�K��ۘ\���T$�)B�|X62��@;���L*�2ҝ߳Q/�,���;��
!�u(��~֛�ڔ/=ME:m!/G� K<�ܲ�j^2���⺘�����!��<(��6zݾ n��0�_ߙ�j�ͩoU��$Hݳ��Z畍�#o��K"�/=Ӻ�+�/:�'�ʵ/�=���-e5� ��*Ȑk%M� �܄���j��᭰�5�Kul�'a��9c_��ء��e�)��r�n6_#vq8��7���l'�eQ+�W�`�RG}9���ߘu4Fc��3b�wf`[e�}=�ר*�����l�6G���%�EQ.�P��C��P�9V�4#N���7:+X��ض��5���e?Q4:�ۣ?`�=���f�``�O���H��#�C��"K��j
�Q�$?`�/�a����ՠ��;f��]+��k��ϗ�=��~G7i��Â�a�L,'�oJ=o�a����Thm�^�[�~S9��}16���o��N�b�#YQe�����C���S"��Ȉ_�}ߎ�9���yR�xtǩ�z�W�j%c3L�ݾ�/�C����
y"]7VC�N�A�/[�Et�;|1��އ&'c1�� ����0��9!H����M�6�9��(�-=�����t���3�|�Y�%��>,�:��Q�,�,;�;:N�<��A���8�G��3D�YTRR�ZP�=�
2(L���OMF7�?HïD5�rMp3���72�li�l^d�z�j*Xl�
��-��rN�V�ᓏ}#����
�򎞚xC@y�:���.X��_��>=3XS�b��=��'@bE�����_���G�wەe.w&�5��0�3A)��ϝ)��NvnW��N��DDE�3�}��,VŨ�طQx��5�����oл�������E�@I5�k|�:1��O7\U""���̫�A���Ӏ{,�����u���c����GNZR�����gY��=�o/��;sd�����\�)n#+�+�{r�0q=K�k+u��=&����IǝT*����{�!4�H"�XQ���>�L?�^���m�"1	M[����D)�����1?l ��)��͝w�n����Q���}R�&���&�� �b�qe���L{�t�Q�T�����E��?l -z%��;������'МTYn5G.|�V�}�!R�;ŉ!���h�\�.8����8�H�52w���A����ک1�I�����vg�a�X�N�˒�;7�L�pih���ձE�s���}�Pѽ�%Q�V=�Bw2%�b*]�[��TܭJ���/�� ڎu;���pӉ��w�E0�zj�`�,P��E�ůX���ѯ�#q�ObB�*=+c3�������E����0���������4>hkF�s�6��G�������g�?��
�ӿ�d꨾L1��)�	�V��.@��opzG���y�˘P�;�K���i1�L\�W[�#mᶑa��'�|�k%V�,e�L��l��lĥ�3VM3�Ă�/2�ė��y[��Ֆn��M��h����AF����$(W�Bܰ|m���nKU�t�� ���O'|�
�u@���eNX����+U���?�/Q^U��lY��0*\����6�>�í@Ϟ|���`�$��Xߟ�C��Q>K�;�u*� <�Y��袙ߡ���U�<5�&�aqt���>&Fz�y���$RʲG�x�9��FJ�:4��o�d`v�	 �>�#�M6��u�^+˩��"b�{�6p^��a�ߞ��i%a<MB'6�ݶd���NGS�4-̲�x�i]�&��=�\�����%�9���O����5-;r!�L�[r�g�w�9�y��>;x"�(�t�eS�C����rvÆ  erH�,�{��%R���h����� ��`�l`�:�e��T|l�����KL��FCz���o��wk��ݚE�Ӗm��It5P~��6G�'���'�:�d6��.�K^.tO�J�~�RtA�,%���>�� �^���=C1��¡���»v�)s��ɠ��5��빲u<g�>��:�����S��܇�|k,��V���Ѣ�&�u���݌�;Owb,u�8�����][8)�7n�&����� Az�~��WOr�����M߷9�ܠ<g���-�:C*����S.zrL��S�P���.&�Pv����9��c"4LJ>����� �j��h|*�8�<0��/{N*�e�M9F�j:�0}�@9-Qg��g]�
�U�GHC�Um佯7�ף-����w��h_T��g�\�ʏ��A�7��ؘ��Z�<�O����xW���w9Oh]+���0���i���]H7�[|p�!k×��]l���/q������y����2��|�N�?ë�`�2D�o8 �o�#�0gE@���>��j���[�;
�^1-�E9�8]�6u�+6�������t!M����@Y"�\���b�[�_�1��,��ЍD���|'�����+�����urwn��.�59�4�Bg�'ֈ�k6� � ��4g����S���	�^Yy��8h-7��W�e&�N��+��<R�T���@�+��U��V�l�P4;�Ȁ�Y��ٶ*�K@�&��og�!�r�~=w�;�j�We#��2Xb<S��6�J�\���f`����5Nn'Z�������z��\���x��N?�1rd�c��Q)
�>t��T`*��7���KbA6\��VI�<�N�C:����2Yg�nv�,���e���$E��q�	m�i�8�J���Y��`�M�va�s�j6�F����{ö��:�KE{���Y�u����Xٞ(^�g���9,����6�̊[�>�����,�BV�[ �����{�<<�T
��S�_T�B�X�W��f	E/3?����J�ű1��Ċ�Fs���중U����0��%sj�.�ya����2j�O:X��ŷ��<Za}�3��[r7��\�h�G[�&e���Gx1��1w��w���9�i�yͻ�'a���:�j	3�����M
u���Ӧɵ`�+w��w��/�M��o�=������v�>�JT]����'ޒ�݉�.6A�m�$R��/D���q��)L��WXeRgi����sA�!��A2o4����������qjX5M���:L�|����Dmݓں���&�	����h�!�P���5#f�����:Y7v��/�pm��rń��D5����>x�('�_	Gc�c~�탉�X��0fI�gR���Gռ5>zlPt�7,JD�t+1\	-Q��Ņ����ł��I[�T���-�6GN&�k�k(�oa��P	OY�}φ%��Tʏ���PZk�}H潌n!穑/���g}��'f6�H�sj�������eC
4㊉ua4��w�[�zZ)۟*�y��ٷ�eP�[(L-3z��pFԝ�tu��/}(_��=�7�!�mf_��kU6��tm�X
�=%�����[��W�r=���xnP��r���Q��h�'���(�%�X���Q$5�XB����-,;���JL\��jk�e]2�Q�'{�x�N���pq��yBa���O�X�:��Qj�������5�c;'P�/��JW���0h#g�]�e�*�u�'�j��n����>4�K�;#}Vc���a8���p?]�/i<�ll-�E��R�W��[�si�V�r����t��Q�����F�nB�=��,���ua_�8���`i5�Y)��{��[���}&˺�1%��P��h���7n��H�)�O( P#�Y�^J��`Z��נ�^����|\H���#���X&�Ff�ߢT(��?���!Dhԝ�N�|�	�*WK|T*��@u��J�Jp����?�u�h��� ��x/�O�(����ƿ�I��5v�"��vc?�3�v=�$� qj��jG��g�^1$�n����e����)2 �D�U�O�?bu3��6�l֝��bF��`��n7���%X�#�>ڱ�����<P�_��E�/ַ\�e��D�A0�;[�U���?�3� �K���y�D��=�6���t�t�d�6ԟl�f�m�']5�������Xv3㏼��Cs�m��m��!�	�EQr���������L����eH{��Fu�(���H�U�w�j|;b�o)���Tn�POr�L�uB�M��H`�--�r!G}��	��hA���hB.~>�  �a�L�4v��۰MH����e��Z[�S���j��dT���1߶�Z`_�wU�'�8y�%�^U���w�Qu��}q(։�R1@v"J�#�Wbi�/$���.�B��2߼"����T���閊�"
C۹ŝ�*�?����9��8��� �7�"+h�$4D���%���s��ȪP�s����n��'�'�]�Zv���O͊����Mf܁��o8�ژ3dk����������^����GH>PM���1���i�y�E~��N������+vΟ�8��[��<Q�wҶ3I$y|�ę�5
��z�����L[,���]:�̪gJp��w�ӇR ��,��b}�r�����L��c$S=�*�둶`��� K�@�`����p��~ZFM<�d�[w/�!������GҀs�EExjWy"=փ�d�i��
�W��m�O�yőh]�o��ɰqm1�{�V��a�S�~^����/Soi�K�H��vz%��bͼ��3z�f-�pt%%*ٷ�� 
h�ی�L��[t�Ga�ng2Jd2J(8����8FO�� �&�g����}�T�$m��Q8M"�;6��66^`��M��E�V;��G�����?�[.<t�!�����m�u����sl4 �"�0|���;��>�v��H�R�]�)r�mF��v�g 5��sd�]�ÿS����G��d�s��쑚�`ₑ t!�q��:TM��m�>���M�9��@�}��ʭ�h�9/6EQ B�I��&��,�b�#d�<!YmH�!����0�
r[	|��F"E٥�(�*k����О���!�i�\�	�ÚL��dp�y�.A�C�I�F�
��_��U~�l���������߉���2�Ғ�ȶ:�[��{7g�6[Wi�,�0;���ė�D�a�,pC�����}6X�;#ʘ��亚ݑ*Q�%ʸV3J�����|9�w��$��|�bH%�XA�|��(�8R�Pj��Rt�ڕV���C�
�4��#ΑA��Nؐ)����A��Y3�0��4�V75����_�P)���j[j�������#�!2�v��.XΊ�t�إ��������rt94���U��>��n�(�o���r��)��8�m��L�kX�d� ���[/}�#(T�Jҕ�@7�ؓ�&�PI�l:.�+F%Yʌy��}ƯI��d���Y�<ٲ$�M�J.]R����JHI��W��
�%�ى��'��Ԯ�t;��}��a�}���*�F�#>�X�&CAՖ΁�a�f`s����Y�|"ih���V��'�h�$gja"��S��#Z�M1�%*�\,zA#�ل���A��� �H�λ9P��)4��"��̩
�zV��9bg�.�{�(���˚D)���Jj�<�w|�.���?��I-۵�Z;�_����x��Yd�ʈ���u�p�RxY�V_!V�$�?Č���uH��c��A�s��=̷ ���p�|*���~���k�0�|G��b�ɝ4��cF���$�(Ӆ���A����~��z�M��<�TkP���q�����րUH@&��&UDH����8��)�Vt��k��[�E7f�W��'�,�2+��%��/Ku[�B�o�ChP�1�������r��5[L�S�V3��m���Y���ž0j���_!�q�_H�>�v�bo)���0龲Z����FW�q�'�Q�V�Y|1�%8�E�����do�I.qݍjW 7�7(��I3ߘ=ʁ��pY�W)�M�k�m���[��O�Gp�":�.S�'�+�d�r^��^u�n�uC�U��/�Ska�����LH��9\���U��Y�J]�����q[�pk�z��.�,Wb����@�8�Sb1#1�g��^*�O��"Ҧ/���(�4����2�J-.��;�j�sJ$�ܹ$��� q�\M.T܆�ド���鑨��~�/�d��"�2�W�↎�çq�J1m�)�//�cB��r``��_@P�	 �� $f
����i�������W#��걇���f��Nɭ��u��S���Hk#���@��_�0ލL���e_���)�������x.�6�l�MM�`k�+ɐ�CAUG��͝	I���J�jhBo҄)12<(e�Q����8rG�����Qp-�����3�V�t<�ۛ��g���-G���0�������VZrB��vt�B��EY��=���e��L�bVQ�>m����[������.��?��*W���'�2?�1Iv����RL��*V�J�N4z�
�_�a�1��Krn��0R��f���?�a�8�N��3�n�{ӯSdI'1>�!y%��:�p�л���Nd)��Z�~M49�#����;�;�$�?_� ��L�g^����ܾ����H`�K���U��������l�?����R紊�����6���W���Evݦ2�GT7���s��G^Ɨ����0,��2��_�[��"S��p'w#K�	C���el�R4���Rb��M�=f�$�,e�8T|[�^��iq���k?�b���tD~��~S�W��Hr¯hN7�/��I��i�:]1���K��޸̰����h}����E�?؀]��+}A���h��bP�u2��u�"G��l	S�^`��,au�X���&Oci�����f*tԶ�>���l��g{��yg��;y�.f��~3��7��Y��}��d���S�Ve�(S�i��>����	��SX�1��o��-Q��"��s���R��}�5>�v]�~�/�t2�F7C�z.G�Fϫ�#��(H0�TZ''|$EX��F[uo��� �/��Qہ�"9����s3��d�;��M9~��n���\����<E��Vp�?�W��Z�2���7�g�1�OZ�>�𚴟��Z�!��$4H$�흿��b�]���E7q��"���(P�g`�)���CoKCSHp�K$�@}����^ڨ����9X�O�/��`I:�հ��*ʐ:����-�XF�d�$o�q��=X�=!Z�7۵;ŷ��=�v�W(թapݴ$i]P3���a���y���a�Uɂ��0�!L��`��:��[p�4�k[f��H΃	�i�4��ߘ\H�O)��/<���S w�ytPB��>��h�Kj�i-�;��T5Ծ�?��Of�a��w���y�F2Xt�Q,�;�Ӷ��Y��4��;��a!ɾeky^b��N�+��:���E2�*ձ9��j'Xp���S{���bwH)���d��[ ��8Ƹd%h#�μf|�%���m%� *��> e��n�����Z%�O���&~�[�N��.Ό���$���v��O�*�r\\�#TѻX�UH�_3����7�_�Φ��"#Z�2�?��e��y�|>�/i�2��8z�2���*���՟/���Ќ��=F�l݋��ҕ�aT�t��������:��ԫ]"�iAʬI�)h�|�քrw����e����7?�Xs]���y���l.��Ƭ��w�b��t_�-�
�Ob��g���bQ��_ӑ�1�,�EQ (Ed�7����<`����];ט�l����)��Y]�v�m�p���s�oŨ��R�ms��P���h���$!�)���m�h@!��������:T�Y̬mM�d(��he'��K��W�
��!�j(19��c	&�h����j��7���}nО{��E=��o�����i�gw��������$�+&ep$�n3'�\���s"�T���6�o@��(��
�$ ��W�g�ڎYӷG�H-!�+�ݺt����%�~M��8�˾��^�5,��$��$t��z(��Is���;y��˕�W�FDE~S(޾E���>)K)L�W���MU=�e�n[�+dW�n�T]#�[4|�v�2[.�i��KL�l/�)�^�4Ǎ�k\�?�4ܮf`��C�����#d�p���o�Q)T�P�S7����n�gC����9fN��e�U+�9�Y�]�Vd%��<�BV�c���"���n�����.y��*��F{o����i�X%��a%��ZW:���K�sh#�"��\?L?�J�%�9.��ڛ���pޙk�]ѩ��N��cؖ>��Z�F�$�{n@4���>�0͞�������-T��4Ă�ذqɮ /J�������S��ؔՌ�"\�6����8����"Y�����K��B{�� ��	��y=J>�%P�y��和Wlk�!��q�9�r/�!A���ɖ�PmIq�循��v6س�6���,�/vc-�����!���	�d��j�d�U�fA0Z��n��6�jn��(�u�͂��� ��߃(1O�k�:�)�z��֪ �Z8q���6R�`?A�$}�n��{ALٚ���d#"^�ۮai?4�v`+]�~�^O�*Rqk���8 )&���O��X�#�ȸ��VԝZ�_�y���fwsߨ�N8��#�l�������0�e-��:��"��vO��o�.W�i�(%��Z���i�/b#�.���	�ྒ�g�~|�k�<�G,�(��s���i��"���̀�c#H�)$��}�TۤȔ{����ɯ�>�c��� C��,J�](S{´~�h��òMTh�=ۥ}N�,cԢ��6����{�rם�H�=#�pJ��N���-��(���Z�˽>�8�Շo-
P$��aI�)-9~���M��"뻱G�����F.vRbCɸ)2����k��
<�����'�,�BJ�H5�|��ވ/m�g�mP�C�Լn,���e᫊��7�9���%h�C{�>�@�:�{_����1˦�:��4��47��B�Nİ�[�W4�������be� N��| zF#�?Q^�L7pp5]����I3dפ��c����W���`q���k>�b��Kj�sS��Y�> H=�9��Î߂��R��-2wtj�v�˪�3� �D��|��y�?�U���mmh�i�q������Q�^j�ifO��'��Q�6�����K�Y�x���(�	�>gFPى��oXr�?�k�;s�u��=�,6h��B8����Q�=S����E	����L��Q��&wn���\���U��5������*����M�Ȗ5杞����ޗtzC��i��\Y(49R��vy�¶�"�F�	b͂�8����a��32�AC���6��_y<����ӌ'p��F8�۶K_�RX[[tu u�;��30��;������ 7�H�%<�#��i-:*�hy@h1!^[T�%�|�<�לXRLwu�pc��,����}��$t�nZ_���hh���kex�9��m�c.�[�i�Y�Zs��8����i䬐�J�YD�b�e����F�Sco��7Ho����*ڭ�|ZK��x�(����p���`1��)�����Vk���;W��h�y)V�b݂U�m��g�?׵��"�W�lX]S�~>�����G��� &�ߞd^��p�9���������Ƒ�E)B&�:L�����Ə1g�Z�������Fr2�"�R�;�y�}�a��es\1�Q6�%�_W.
y*�~�$��e��Ʒ>��>Ǔ��49�r41�VZ���� Φ��Ħ W�i5��Xä�z���z�?�J�sO���oW��T��"_C��bf�@ d��5�9<�����G�F'���=��쥛������b�޺�>J���|N���G�f���_ߋqL�3v�-^G���6aD'����Wjj�i��C�)�%!����>����o<����7�����g�B��ב�������a�a�}����[�7�%�(��xzڃE�z�n|�PE���I�E<G�w�OMď����!|^�W���\��*iDes~����CÒ�^�
_lݱ�<UG'*FG)*�!i�@��m$�x��i� ���b�J鄴��e�;Kԡ�ϧ;l`�r�ƛ��[�
r^YZ=27���V�:o0�=(L�S�g��ImO�}8����/�B*�"�$'��!����2�$/���Q�3�)n�/��!�,�6��А�Ę�����ҍc��C�	�*jtZ9��W���#�D����N����,���I�ǌx�����R�!-
����N7������8�)k���w��p��=l�*q�[�|�?�g���\n�}|f��'��h�"�4����Ϋ ���kT� �R���~�`��.�:$�a�>�I]�~����6�-,v�I��%�$�\Ķ�"��~㿞�b��"���� F�?!��z"� iyVONy@}�;�����C�N�%z�a�(O�i}.YX#g�L>�B�hS	��1� δ�2��Q�mĕEbpϑYzes:�H�;��\���Y"�1���P�3�Y��S��{-x�r}!g�(�q�<���	c-�U�H���M�S3�2��$c�XE��A�@�{�6�ǹW^��-U�B��)��2F�%b��.2G���t	#��KF#�5��h����i��b�a�c�n]18F��.��^��ސ�J��p�6���'�����9L ��Ϝ�S��u��Qg��d�`��Y�K�U�u]|�H�K�G��+OӪXxf������t�P�$hN�����%a�z�]P=]GPJ�@���to`r	�����ib�49�-ݠ���`����-�s �%�T����=f��6ɃPf͞(�!��5(�q�8�e����:d�J8Ɔ��FI1q?����#�G�Q�D���AHޮ��EzJ�V�@�XR9jq	#MF:2���:���@�Y]�ʝ�w�g���BT�$�&�2�ǰ�v�f�mK�(τ�#���w�y��B�H�C?���lR٭\{7i�%챟S#��&��z&�%$���Ñ��D\
�Y���!|�bd���@��ā87-����s�1\!)��{�]~��X���ļ
Frc���yT<�o����՞�%H�jUo�@#�<ߙ�Đ��@<��Fn�Z�.���#�`W٪�)�ub ��r%S�vR[��X<:�.K�4�� ���݂��U�����M@��*��O��Ru[�7/����q<&�u�!����Yw�*��B�WKCs�J��qu��k�l{�1�؄� s�Dr[�x�������Nك$^ɇ�l�*����Cd��sRX	"�?��W�}ٌ�zX�+47�5�l�kyl����X`{kZBr�S������
0��vTC��i���	<Bݺ�ۅ�o��B��YB���>	ᖆ�_�'I��>�a�Zq�]��NqT�\��}(|v�]FwĚoPtB+��V*�D��\cN�� � ��h��I��\Si�f��D���(�ѱ��آ\�&∍B��jk��������x�sD	�qW��;�Bj-:���A��e�4�F��m.Y���3z�)���[o)u��x�i`�5�R0���y���g/<g�;��,�ZP^��Ҁ������{���eD��R�*��J�1�Ue@��[�+֡��[�(�؂{A��/�ͩI��X)a���q^I����"[���u�L�:�ث��:���0�"-t~�kO���
>���L:nJL�̽m��Ti���*h����S�u������h!��߳�Nx�`��-�����K�`InR��r��۞����2g��Ta9��8�����>!%?��t����]Q���V*�	�C�屎BJ4��C��ɰ0��}s��xU�f@X�R�Θ�����y��p[C۫%(��A&�Fl(̣�JU;�Q��n˻��E�0K�	������)����4t�`J����[�PE���5yq�圞�
��@<q]�oȠ��<3=�4�k��у`_c������R���J��^�� /�_k�#'�(b�_lبՌ�e��a���uc(peS1��9_G�%/�t1����#�^�S�X^����[��k���K��hܥ@Ί��#(lD���1����?�M>�\`��ˤ,Ş�P�D����ݫ�+���RCk�J���r�
Q����KmOt�ǻ��Y$p��B`��+�;�� kKUI�z�z�Uw-��SL�"
y�+�9���9<U#C,+6������@Q�"�]�fMI$>Kޕ���Z��s�oѦTcD��8�|S��ux�Aec�ۓ٤4Q&���B=�%����OHc�JV���)���[� �C�_-f �|��C�
��G����4��bAq�h�5���yF�K�k�K��L��� ����G��Q�
�;��	I��2XG��s��V'�{����P$wl��S�M�S>C����儓�2H�)� �E��./����e�"f{ڤM9�q�	�m���+K49�;��*ײ��s|܍N$�U�3%�!�hQ��8�%M��l�Odn`��
C>h���`S$ۅ���Һ���C��(�Xd�C`R����o�G�,�G�R�뢾ʖv�]YC��z����ƃK�GO��٩@#H9��b��<�W3a@cߙ����U�,�x�d�g��Y:���L�
Y���lX���Ɍ�&�r�G��@��+�8��[����'�6��̔�0U�{^l���`Uh@���~�ڧ�]�0O'��F�bT݊�p�$�Y�P��9�I.G�����dt���A�\� w��K��&2m�@VcT�����@����v��l��`Kp����F)��8j��㖐cA�Ȫ�U��d#���;L�<WOTc#9���V�0����!��X���XҋJ��Ox�J9<O&N��%��ʯW��
�q��V{%�B�*rc�U�����,�J�ӆ�A���#E֔���Fˍ^q�sǅ�^\G3_��iZ|��Xot���2j ��:�6on���|m��R��%�A�C� #.Y�;h�S�Wűm��|��EJ�0=���ݶ�����]�n��i\ѱ[��b�D��ȅ��HSg������Z���zEQ�[*�x�c�2�� "�˖�P���X������#��"��
�/���p��<N���q`��r���o�*���.��g��j���,ڨ��yl�[�[ybE��p�H?��薦,�����]�����c\�6�[!#	������9)ud�Fa���b������J��{��Ff�5�Q��)�n�g�Hn?qV���5A��A�s���CU�ړw�S���a����!�Z�9b9�	/P��Ѹ��O�`�"j�9�m`_N�f��è�l�P�!��B&*�.b����p��Yw"p��������*,χ��^}E�}���oOr��	DP�f-5���O�z�l�=�CE���F��8�x�z �EU�iF��s-��u�5���M.��Jsw����|�.�r�ct�Ra���)�f�.����8�x�������~mu���|CHȁ���np��y�	�]ϯ����͕��ƃ E����R�'8�wo�P�OmǪ����C���� r1���zd5���P���l׬��1(2���eȃ���_^�͞����%���2S����*`>`XA2�A�-+��g���S.<X7'14�A��B���<u�@4<z�����,��وm��V��&n34�p�
�t�����b��__�2@R�.���%���~1X��XZh��2/�(D]mE^X}�R��0�<�6����_��Nk�{��K$ጌc��=��p�f�Rݳ���{��q��y܇�<��\�b��n�'����j�9w/�Tk~@��;M>�I���j�_4�tZ�tP�}$P(x��o�zY�@�,��ԯ��k�c��Cv�G��6*��[���bi�Awm�� ��z�	E��)�����Ŋ)��ѐ]dӧ`��#^B����R�:�`��+�@��u��у�����2�d���7r�5���=��>84�O^�D���'yx�*S3�&^��9�c��Ǆ����J%��] G��Y�©ve����<��m���~�(����u.��t��K���>�C�X����%3�TK/	��Ed��h�<�|g��^��,.��uL2��U��@��1����5��etG?Yn��mJ.�?�+ω�~�K�T1�R+���H
��+���ji���׋I_l�����(���	x^�.��*�Ǧ,`�r���=F3sxΥF�eLzj��O�R{����-J��W�t���y]�ʙ��Vo��hV���I�5~5%k2�Ǔ�q��Qg�B�ק�}��@�>/ ����'�r���G��,HUb��X&���L�{~�f⧇�^�g:^?w����ʛ�K�4]p���n	?�ե^i˩��Peo{�e�s]������w���h�P(��mǧ{��@����g?{�ꬸ^�"'�t-������.��|v�hڿ�L�,d�coQ��3�̵>��4�0����22B�k���F�䰏D^`u:E��s����+S]g�5���΅��>n�ޔ��{�~e:.ϗ�P'���vJ3%��P�],��.����q��a>��Np�;qh��(��֒�pѼ<�PՓ�r�L0[�/p}���ſ��9�M�+�f�T���&T�髂s>��=��^�0W6r�E\�I��c Eq�I�)�'�zRi#�[��MP��W	_V)�lZ��d���wֶ_7R_z4�t�������E���
�ziQdVC�h�.�2ngP~=���5H"�N��s�7�Ř��54�ܩ�#;��M�W����ϵ�.k�pn�-��ݹ1`|��{:��eHf��Ёk5��}HL���)�ώ���EiD76-��f}@#ݑ7�&��+}�=XKU'�H�K!���^�`f����M���u��ؚy3����cX��4Pe��C�H"e��"�����ܰ=
����m�tW����(�x���
���m��[�:-kYC���7r�,D�j�����4L��R[�6�1-D=�+}�`A0V�s��J�&Œ�Ã�+�q?�ު�����o��λbB=�k�pu����u�����'�Y+Z��)��,�I�'ԍ4\�퇾hc�f� �@���@Е�,�7���-T�oŕT�A1Q��}[WN�}aD9b6�	XmR�1��7�|x�~�B��K�V�Q����x%X�X*A�K}vQq���f���YW��|�A�
4oe�}�yO�,8�+�Q��(��O�|,`��Z�F �C�(�do
�j�co�xU�)*�~�T��5\�%|V'$q���Q���v.��MS���8'�h߹f��a_9�� � VN�˚6H���G��J�}|A����A�.���CwK����"��[��j'}!�F��V
3�OT�������T� '��l���>=GB�K�9���P��Z���@�+��: ��Rp��Q�͟��B���n��q�h���酘�x�+;,���P%�z5֙�#�ρ0]_����x���"�M$2�]*x|
�2�i�}�2d�t�)�AhG{�ϯ䏽��� ��G��CJc�unmGg��$cn�D�W�����y���:�=���X��N+X��=�(�q�O�/���;�w+��:1�>�p�u�Մ��k]�a
FT�͓U$����OBu��⚢��-a)vS���C�UlV1��=�Tsӓ@Z|��v0^�+ ��F���@����}��س(S1�20£�	�	������O3���"��_�ȗ�@{@�!�WMt��Su��S/B?�-SL�QyD��z�}��"�-�kqry��d_Հ������
B0Cr�8�e��x��E�<X�p��JU��e�9����(}��@�(��*~�X3.��ښ<�01H�u5����H�vRL=�ۤl��GL�^�ߔ
j\�#5��GW��>��X�����e��23Ѥ"��*綂mH���c�c�N��	S#�������%�[{�ID�l4i�+;���_�sJ��6)�P��i���� eŠQlt�V���k6�M����\���!\�S!XH�Jv�Ͼ�^��ᤞ�P�0"�aݰ���O)��J�h��W�	��4�T�<�Ftm�`sF�Rs0셵Q�ak&��g{ щ��
�;M�ܾ�O�L��D��>z�X3'�����P����^�j=�ъ˭���C�4Ҷ(��(�$�I��%��K`g����L��j_W8�6��cȮ�I�]Z��>�yl�<����sg����$�d��x��jw��?ւ4W�u����{��7�}�P1�)��O�Ն����X�U������p�})�������s7��=��˼|}�����'��n�򐅵x�&��"�^�M@{���ad�RP���r|Z9BVwV�!ko��`ʭ4����酥��jrƺS����MF��}���Ԗ�;���@k���8a�\:���O�u�dF�� b�k6YM=�Si�.ٷ�ȹ��.��vL1��I�O��e�|��'�U_��K�8@�9c��K�;1k);�vQ}?���P�*�������I]}m���~\;�5�����E�T��{-���Mc��ym�7�(����'�*���&�9�9��"�<�`J�������؂�l%�ip�L6]��@2!��2��&�ʇ��)�op��T>]6��`��������xDƍٿ�Nk���Σ�iCji
9i�m��e%e4��B�ɼ��~|7�*RCN�8�~��߻���Ӵ��}�\��V��Cƣ��Z�ٮ�����`^K���#f佡���c�^�
���y	l���i�� ���ۜ���	�^�.o6N5��q���<��,{*`��z�?q:�C�U�Y�9�@�V��[�����s�j��!�%��S	��	AF�U%^��r����^�CS��L�/'�d�{k����h�z\u�ճ\�p�^<�1NyJ����tъ(��>�����@����c���5\UޣCM�i7��~(ǩrI�|�1��4��r���v�{A��ߴ-��#�����cݍ�=�kM�$�$�y|��D\i���xa��/!`��/5����m[Ƃ;V:��7�>s���/2��&!ٷ�c*b�O��x��@Ȝ��O�~W���eIٲ�;�30`�q��=���8iX�b{q�/[; ۫���D�w�m�~�'Ka^HO�����[zV�l�KӉ���ф��J��Gڮ�@�y�؅R+γ�����MX�����WSg8�(��^|(G�. /��|W��B����_��o������XV��|u �2���������/쎫����J�v�9�l��x��Q�n�i^Te(���/{�n�3rv��Y�c�����+/��WhX��O�W���)_��h*�?�!�{~�E�G� ��j�4��%J.�GG�h�&sz��׽�y+���YQ�it�?={%R_���|���"��H��s�^.�@0��rODƉ�B�/�,%�J���������X��ƭd#T�������H bV��oi�oGI_�P��6��4E�ڬ��E8�k���=�~��_��-1�o��5���-$r²��;�웭�!
`��k�l50����x�Wl�!�6z����
�ymi,cm�ϗ��������������#{�_�|�$�!�7C�t
��PʺF9���:�Z]AU��+��{� �W�ii�� j�+����"z��Rdr����=�h�Pebp2C��e=oO��a�
m�g�'�+#D�&�2�d�!3�-Q��k�20��"S�3��V���j�J�y��8�K*(�f�?��O`e�z�gY�as6h�@LPz������E)d3��'�������-�*z�V��W�ů��{�f� �\�z��`���x��4>�H��X�+���np��L��K�f���' �^1�oE迄Ggpq}yf�;P;\H�L6�x6�ѥF��aB�dj�x�K��~T����z�v*5t3FAChW}S2V����54
����n嬊A��4|�y��ݐ۠{��tF��dJԕC�}6�nR��J��vr�]������*h��)!?�#�$�+� ���,j
H00-֫[�K ��5'����{�7䅚�Qqb��}mᥕ�����>����g���	��5��LR�e'�Tb"�J��,��ݥ�,�KLQ�Zn��-�6&6�`��Kv��m�ϔ20'�LQ�)(�u������4��݌.�G�x��u{��6��`a�X3�x�T�g+h�;K��1�2|�D�K���#F�Wp������e�e�"�	��`����۪�hDcJ�8^��K��T�pI�3R,�����շ��r}bC��h��K�E���Fu�iHGϕ%�7@��V�N*��19����/����~�̀��#�^ԩ�B='v�¬�"����Y%
�󠡉��{�Th�[:�?>�8�A*�G[����k�t@�����OZ�3����^7��D��W��ֶ��66)o�Q�k_��9M�u�F�����,�Z�^�?A�Z_�U��5lJ}Γ�2 ���XW�;���M ~Ŏ�����H0v�1�s���� �σ.X����W8~�����6���������2m���a��Ӛ<���R��J�͜�$� ����<���$�Dz���uaM�W}x!�Vc���v%�v���yW�?m;���`�X��G��������8�V���r�7�����U�gfq7a��!;Ӈ4"a�Z��
����u4W�HB�ToWG�g��/��nOԀ
BD�7���3�S	w�cGHM8W�5�YU������ݰ<�i��2G�۫��`) O� �fe?�
,J�#�_V�o2�c�=L��I�:U���������͍k۷�p�������f"��*�FTv]�&+ �dEwu�@t��Un$�\s�>�T���t���}�ިQ��_�<x����q�Z�d�u:��-�x�C��~^?(��Q���WV3<���q�m�����5������KO��>�<�=��ұ��~c�������L%�*�/���'C��z�(Km�����d$��.��,��ggQ���?�N�w�s�f�oO���iO�\9=��f� >�2s+�߿�������.l6��G茣2텺��{\}�ϯ<i�{D�&[���g9Ё��$�=�!_�ݑ��&jX+�σ]ű�]3��|z@��EblC�� � pgJ�{�W�o���+�W3���]6[�Z�@M���`~�t(��A�p�a�+Z�������I&Tү�"Oz��g�|�{S=T�j��x��y�����}fHo7;����-&;��q	~f�����f�9��D��hZ��ob�)��+��9b��&H�'�h6��K����m����`y��ѩ�z��y��߿��ȹ��qN�|;�K�q�.�E�=��,�a�3��?B@�
��n�8ퟝ�9�����r*^6. s4l�^��jU�)���Pb��z˵P�ę}{� ���i
�(:�եp�k;};&� �0�a:�hK�:�c�ڜ]N�&�^��=4�'�?�D�w�EB�|I���UBwKD��Ŭ�{V	��b�����9�!����W9m�ΦS��h�)t����	��\�-���OT����}�S	�y�Y�=��-��h#X�g$�xˮ-��c#�D5���"c?�+�G��g��\�����Y$�������)q� ޘA�7S�ф�1~?W�.�j���=婔�c���:���y�=�P�]z���=q�D!/�쩅����2'X��Z�C�u
Kf9��[��JJ�}�v���s�����w�%T��(r�q4񻱪��l��_�y�J�v�q5@���b������2<-�A^
u��6�_Xҡ'���oq>lr�2笡_�6��޾z�.���M�!�̹��)�O�5y8��!너�u�1_hs���&�q��}�_麼���"�<<��q��55�� ����W�wlT4X���ad���x+�*��!���z�f���s�`�'���=+x�ye��p��GON��r��m��S`-h""�{��bS,1�Q�/Y�{�sF��	�VOQ�������: �$�`e���=�%K�F1�!{�N��Y��T�����ߺ=�S|n�:�� o�<G~�t�7���(a�ϓ]p���4���N���=�+>�Ō���<i���� 7Ep�Z��ƐhT�����/��u��%������_Y��*��HZ`8m�D�IyV���������'�BN��/adۑ
O���N�Q���v��浱)�:�t$*R.j�c��~֫ӂ��ۢD����!n�+ә��I||�D�o�����7��o��s��gp�%�n>��gP�\�X�'L�#�/��km2��*��y�ꞯ�u�[,�@דX��4�q-|���*ؑU��J�ʚ�V�~Ƕ�mp�T좮d����q>������b(f_L:�U��2)ƃ�O��|��1�� _��f����������)�3�;"�½�YS英@�v�y�d�[���ҟ�[�L1�
;��a��g�Ҷӗ�G��}����γ��N5��_�4wb����%�8��X���}rڅ�Z�^�؁���L#8�����W=5�
q����?��=�GxR�|5aKN�:S�˼
%��@� �^RN���v�T/ss)�{-����ى
�QA�F�~���ob!��Ķ5I< ����7`$�fs�3i�$�h���-�Y�L�ߩ�i�)��3%夨�]G�e�hːk��q^M�@�&>���Lմ$�Ov6I⑇��b�̞~%�i��N9�XF�Y�5�N1nBv����E-�ha���1`�%eG�)'>��,��pat��Xb	��W��l��X��}�8��8Y%}D�<��_2���|$�k��w�z ſE��"4Uc��	F룶
�ׁ�0�ɍ{AResT�+!����|����[��� S���a��M�ұ���:c�[�c��rŻb��n��{h��9�@�ϫEz'������Z5뛇�^�'>U6�CY{)��mIC�<�KMֲ�WZ��P�x����2�j�����jh �-�D���<6o�Kc�-�V��#�^�l���|1POkf�0���Y��4:��r4�%`DGm��`�B��H�BVY]oƫD�a�f�b"��Of���-ϠG*�?��J0PS�dy
Rw�+,�
�R��̜�M!q��rmPլ�3J. ������W��-	���&c�� -b0�l��y�&Y������ĭ ���p4'����b��B*2����4�?R���S-����V�ktbxu�����X<���W�;�u�˧�﬒���}�֨�+���t�&�w*m:׉��K������r�������d�2��S���uUr02�FAdk7�,&֕�ʼ|ԙ#�4�/��Y4K�t򇅔�&vq#F��*���\�u�J��p`XA��Q$E\�l!(wih@<Ѯ�,fal�p��B�VU�{uf���j����]N��k�D��͌��cN�����>�?��L�ȁ����Fg��B�M�\۷V�A�[�e���7}p�^�~m��.9�c&(���E�Ef^x���QfnC/�m��Qz�l�gW��.7僐c�)�F���Ahz��É���������H<\Jc|M��5V�
(:d����y�g���T�V�#є�vV���(�(���e�X2e.#&zМo��6=�󠳉6�p�X���}*�ElB�8	yӬ�V#oNz�q��9�C��y�6G���E**���??c3�U �h!Z��j�J�xu��Q/�����X�e���3U�`f�H�H�ԧ����0=o�����ﲠ�����v�ɂ|�e�5��ǖ(�CPF�WN�@澵Y���TK=l�H��I�F���q=ڨ�X�e;��¼V}�i��jzw��Ȟ�m?�[�0�*�Z��<juK*׽��s��{S~!$J>{�0��g�����7'�*��0ty\إ��$�D�V�"�KC���p��m�L� �Hm��᤬y4]VrI?S�jr�,e��낚J�����*
�BWLrI����~�/:g�W���/���IB�������s~^lL�@���+�.�'�{��ґ���玼`����;��9�φO�-��ηK�+�Ƣs����S�9�����{\�O��^K��#٤[�1�ӑ�$q�y�����\��� F_�4��*r��A[#���dw�
��5����y�A	�Z,6��[��ao�V�*#��5�t��p9�R�#��b��V���
n�*X0���~���OI���a}HIH�F��4hD��g�7�:�]�"G�
�hw�hf�m����X�����0]>���C4�k�l#."Z�/[G�)~0̪�vs��b�N�A, �D\1z���[�U����j��\n����$ێ	���dk á.�N���]J�_�?���w2��u�S��,t;>�v�!���R�]���������檄�圫���_�s��RS��3b� c�� }�Wٹm�ҡ�?�/���k��aGGǊ

��RF��VL��,����^�t"����s����<1�^�,e���@Eƻ8����������G�h:+���/�@\��k�z[F�M�����묐�ǟ�����)�����	s�|X��J��8�Q��ĜC� �]�I�+7��0�GI�����H9��C"lx���S�k�H�T��]��G�����w�*eh��ۚ/�O].e,9��D���'hD���/Éx��c��v��l-�*�t�X�<��~ђ]HW5�޺������6T��)ۏ+ϛ�A�n8�C��<�k��v�(���k�t5qb$+��^
	m��w��`.+ɴ��泅ۯ�'��m)�pA�[K�D[�͂��^��N����w�$���q�x;�n�ġ�ѵ>I}W������Y��5�9�餭�C('aR�<֊&����P�q|��>�m��ڗ�V�y��Y��J^ov E���.w�u��_�U�8K�H�F�Q �z*��T.����W���r[8F,�lD~IAKp6�n �-��M��a֓��%w�;�:98A��0���W$!U�>��*p�Ar���P,��2������z���hA�i�Q�ǚtDd�*�����Z��y�c
���X�@xOp���"H��3望��+!#�L�C6E@ }���/}:��:K1H�qO��u�\c{*Ұ�n����8g���8V{pde0lE$��{��hiĒ�`���|�jY��\���\�_��YP�[´[xfx�8g�׊w��qѠ����9Qs'�U`��_x������eJh޽����TunF�����%Q�a�ŋ�6���sH�����7D��~�Y�&�!�����OF`�B�I�;��;�2��[�I'�uU��x4�Cq@!x$��ű�:.��F��?��]��(*u#��3�o���m���rM|�}�=�3�yw[�<���K���ض�[k�>$��g�_?e�p�<~�7H���������u�����g��e�p^қ8��遹�5C^��W+�PgW�<$�f�f���H��F[TVt�=�E�S1���ш�x��R�M�ݺӫ"���Tzi���<m���,����Om�gG��9~ǝȠ��o�a؏��
��@�Q�1��f*OՎ����+a��+J����E���̓�,�e,1)��P�x����v0�ݨ���@="PH,tI����WZc5��H7OȬ�/~}탞v1�l��Ҋ]�)U�I��mnErW���V�j��Tڭ���l�fQ2;����8�#{Uǿe�*�C�sUS$M[��N��tF�[�:���\�ڤ'Ҷ��g8�[���dK"�X��q�L���+ g/l�n�4���̷�T��M�o��Ğ��漷�r-�O�|hx�{=�T02�x�vf�c����Dr�޾I��)�g{D;@����عW�}��^�JL��P�{�<��]O;;�bh����F�{xT ���@�)4�Z�+?fΕ	��k�L����y;ڔ#X�|S��>�:B�/K��]!ٜ�|)8L����m��i������i]�[���}o�6KK�c�.F_�.)�iU���i2�C�sW|~��C[��=��� *�g:��{�ٛ�H��rI�-��.�Na�δUHs�uv{� ��*F\РˀR�T=��<�hL�N�#d���A��i�<�HS�QY]��� ��
��c ��sy��[��i� �r��*��[���lAb�P�L��P���w_�'�ؾ��!��GcIV0D:��������X|��-����cd��V#��^�V�F��E�Ъ�^��[�HG3������LK�C���H3��-"���6�'l�C��t�jg��(/��y.�@�W��q��� @�.B����¿^c���,�����%G�MH���!�f��1���[X�NT�v��𯬂0
^��Ԙ����U�@�L~Y�m_��~Z2^��˶� �~b�� ��M_�S�nս�`�p�j��U�Pa���i�����'�Y��5_<��>�<�[��6JV�I�ڥ���>�� 2P6����w�?��JL���}O966j��w�P��ߑ���B�s\}C+���M�\Z�;+����Cv�y�f.�U�_3�0�mU[�t�(��������6��$��,�W�^��HJ�{f�ɕN��yz���3e0�N0����U���r��.�8�i�!&��4�A�_'�<��K�(~X�9k2���_5T���b�(E*���,{
$ڳ����	㙀(l��d;�/��,	Qt����$+���U����G<�Q�J�r����o�t�y�I_��J�?N��7���/�%�}�^q���]a?�� q�I�3#x�,�|~�&�l�n�P� �C���&_b�G��V�z��4|��V ��|:���۰��w����E��H\� O}��
�s"{�Z�h38%�*$)W���9��K�����y1#.�M�f��gț\�x��XX~J)��E���������^3�>D�~'����'w�o�����8��)�T||�fa�:�-dpZ��{'q�#d��t�̴۟�v�����K'?t<�U�KM��%�AAА�%������r��D�t?
nta&K�	g��]��6l�²�M���6}�7���*�_�����{�g�#�O�юM�CskH�$'*W�@ulMx�cf#��9_D�k����A���2���SV5��F��c� ���J_r��\��㓅~zr����_����]Ȳ[���?��Բ]��_��1I��~��m��} ��M�	����CK*8�.��>6a����	d����f�j�V�$S$���F6�J����������s���	���y�܏H2��&+���|�܈�3�LC��C���y0�O�4>�{(W6��I��c3��%(j�X�d�����e����ߺ�P���Q���2��_aX�?�����s�OI��qA�8ш�E��X6l�	:�4DI���d6�п5���t��րJ��|]m:M���]�6�*�P!��A^h���&�*�����bi~rYg}~!6�+�U0������{�,�dd�tE{��$X�ltG.�k�j��n
$�b녤�T�ul=����^,=:�
�po ��O���~vPQ6%����&�~Mۻ��� �.FE��:u.�b�Y�V�3��zOhS�YW2g��	��yCa���	�~��eN�PqַOSs82���ڤ�{�kIϩ�!�_�$� �Í���^b1Z�21jG��Z��K��(��˝�isf�.�W���2��D����9���(����s�=/ݑ�
I��3�ې�v��2SM��J�j���������_h
��J�l���(�7����6���<ǻ��0`����P�b'�^��:�+��cx��-�C�ڸ��U{�_��y�9�n�V �e;5֟�p�я_�N��>����J� .w`��7���Yr�g��V)rV�Q��B��q�Ԧ҇Y�Y�k. 	H8�]�.��P�%uz\��F�Y��y%DT���2�L�V�=b�,���f���5�7ED�5|�>#��Uf��*�V�8�a��VU76�Ѯ "�7�^=6]�w�D�]���>�i��v�
���oИ+�m�{Ax�g�]�%[�E�XI bh��V��ڏ��oʢ�{ݘ��x����3�&>�xĕ����7f1n%���-2n$M� �ᶲ�_��c^E���si,K��Л����ifx���Qj y�&5�.�X���dM��R3��˕�?!p��6Φ��3��:n2�%ws	���e7����V�z�d2�e�t{���aP_�FZnz0!�w	a��e&=W�Թz*��KL}�� �^7t�Z�5�&��c �$J�ݰ>/lD�W�ѕ^|i87�x�_ޥTCXd/���\5���W�⾱����E� �=׌-��L�Ѡ�eIsIN�լ�@w˒+t�/�n��cѲ'z�a��,�ֆ���k�p�2`_�*������$�$�h�+�m&E��b|�����������A�K�>Z���H��}�����1O}jE�?_����EVɕt7,���C7G�mvr����pV">����j�4u(.��8pD��/�~�������1��W_�*�Y&C��P�P�G�����$R��u���9���6�~M/����cx����ήB�]y��4t-��dd�"]���}{��������NX�F����Q�/�R'�v�P�R��!�.�V�@�l�&��S��%m�5JI�߇�Ptv)�pO��F�E����'p	�( ��=W�z�l��mU䮐-����0����U�.�%�h�3��9�f�S��F�����P�R�2��Ϙp���5�*�����hhg��k�H����,Z� 8*u���~u����%�]�9������QS�9c[q�m}HB��24Af��c'���acE� �"�����F�`6!?�4��"6�Εv�K�Å~��i�۽}֩��-�X�>I��
C���Q����&b� S��!;��愊�V��g����܇\��+�Z���a�aXn�'@-��*�ѡ�#ub���Ϭ�0���(���wW	���.{��� �OX�G\<C� ,��Y8t���נ��bC+|4*�s�S�I�q"�K ��KK�#U��l�I ��b7�gd��>�<�*�����D�uS�+�*�)���5T�F���ګ��V�kQ�)���{����%T:6n���O\V��w�<v�>�VT]�����$�݉�GV����-m'�Tt	F��l��W~B�0x�_��Fg
<jD��[q�nE���J��ʌ��UQP��/Ne@���λ�<�X��V��q��8�������u���5
;���6���(Z�?#�	'��N�t�)i>�+������x� &zX�	�h�u}��Z�%1�nqM���x����ŷ�D0z�Ӌ�BG��22�6�R��uӖ�Y��[P��v������񟶗Z�ɪ��y9vf��ٺM���K��3��	U~�Rm1�����i�����ٽ�i��!��5�ƫ����L:��M�T,�I�eG˳���o�}���l�{e���@Y���ҝ3f䞽���vn��D�sX²��8m�vܛ�dfŃ��D��� .ˊ����W�s�Ծ�y>�Xֈ�-C�k�>��%X|V�dx�dzѧh�P%��*�<vks�$�_i2IUk�@Lo�����.j��l���@��^�j#��`xF̝R͈�ޥF1*������d=;�U�+gI���dw���)F;dŰ���E����T6��M��Υ0���.�we�c�@���ID��o�
Rˏ}��d����9�὾�
�`j��s���}��=�eSǤ#�������L�1$�"�Rw���`R���x>���+�<��ؼm�@Ei6K8�Ō:��	�o9N{-)�Ƨ$�::h��:�QMpOb*�]".�������V����s��SB��Ĳ�T��O�)�Lp��uɈ��wT�SтZR<\���mM������5��[ �F�s1h�?�	��!�/(Y(�X�듃��=�.���\��'P�íg~2������#�P���Oz0����e��Fw�`Ș9��0P����:��K��	ƒ�|v��jժ��ėJ�g��	�TSa�G��'� R�C���Ki�[��D?E��[��t�Au����D(q�z����+Us��ܗ#ַ����o�>
Sf�uo�p�xep�ꗄ�cK�#Ɇ �h7So21�sX��kJ�{��a�s�E�^�0�׉������X�oEZW��=,���r������)�O�+[�ǃݽBK��zTo������5Kc��x��6t�G����L}�Cr�-�o�hp�7���
�� K<S�ǫ����	7�5��Y�HB䷖�Z���_�d_�_��w�Qy����یct��뽛b���z��y�GR�=��4�t-7�X�����猼��w��/������_��U��8G�h�C݂�[�a~}��3�K޺���weCX���k�����xFk%�QY�ǻ�p@��0/�2�h�R��E>�O$7P��&P#X��ۇ�X����;��j�$���<9��E�m�;tX�$O�-���<�nd���IYil�v�\ե.+0S�؍���Q�0\}(:�k�0\ �C����!�qePT��>Z�e&*v��S�d��K�c�n�2~�)<d$^�T�ǐb9���2�i�v��K�%o����*��D��-�H���Œ�Q+�N`3L�w���B�k.,K�t�!�Q����!�f�˥�-��/�hf#^�a�Y��9L��<\nh� 
e�h .U�R�(���\�e-�7��⇄ߠ|X �Ǜ�<��=A������MϮY�>#c�,�0T���_Yi#$}J���D�o�<Z�7hʽ�
z�
���Y^W�6
=��;�O��_�}p�O���8�}�w2��:
iP�X0��ǐ;�%��Dt-�3���{G�wO�	 �&(��=kP}U/1�z�D�����;��1M����y%�_Eިkgw�F�a:�^���|���ٛ�,�;�S+qm�?H�G� �������S�u�.=����S�C룮1���w�2�k��CX
<*.��"��	G��Ѓ�L�{îʫ�q�l��F����㧌��yU�����s�,b�2��+s$x��}Cj��F칍4ǹ�T��c��I-}!�V�.grF��7�˒���q�*������?~wɹ���f��(�P��&��ͲjR��Z:OABm��X �}�M�d��;$w�҅5Z	ҝ��4S�v~ᇛ+���!e��S��[/;��\��K8�$Gc�{h(��P((��~EOs�㒤1����\���� <R�Ɗ!N�;�_���A57仯�_��E!�I�v�[���A�o�N���)>6�#˷E3�]��]{y���3�R	���ӏ&CV;M�U��8�:�W���=q�l,d�]-WL�^��8�W��.L!GwXx��� �Ё��͠�Cs�t�����Ǚ��K�ߖy��Z6���e�1���b�@:=��6񜄜OO�3
� #$����$��|6�9��܂zi)�(G�Q��u�4�A� xN+x>��.�į��z`���>�ގBd*���e�Z��(_�JRʼ�}����{]��n���x��L�o���fF��<��J�3�y��̃���U1g3�-�-!���!���lw�ƈ�CE�^�,K?um�W#Yx����j/#�9�������X�[r�Ĝ�u�ES��DXq��VǪT���[l�)�]ZEh��*o�1��OJ�٬9 #����@0RdLȽ�2�%=�EB����F�H���ރ�dn7�WH�.&s�)�fV��i���X�f���?�9�2�o�{��]d�y����8IXW�W
c��W|�4�jf��#��	�?Pm��\^�2L�w��y~�=Vš�7�R��7)�^���/6uHJ�l�A���WqiP������[�U"A�ь3C$�I�(^و�I�;���u�>�9O@Zb��Үy�?��e>���t҈��:�;���k���q�Ga��p;�j,OB�V0����A����Q�����$$�j�Ր�:�~E�㗬�gƯ�jqQ��f�cҥZ{�~uwe��Ǭ�E���	V��7(@�S��$��<��F�ږ�)=�p�~	T�����'�c��J����:��ȏ�� "ާm^���z_u7�ح���=���u2E��҃�O�9X�3q}��<�M;�	�j���7);�/�աS��U���MXp���?�L�tj��� ;���?�r	%��c�*6��*�np�<F�#J���-�#G9�@��&�Z
�����ez�v�M��E��j�E��'�GZ⬐�DH���Y�=L&<làOq��H��`ىd^�g����l�]������a��v�B��&��|e F��]-��k���T�)H�j�
���O�rձ��i��f'#��Ӱ�i�穎�+�,=���VHH%4M���'5Iς��mХ����ldF�-i]�ë8�(.��~���(2������o��~�l����3ƪ�Y�9��	���Σ�K��$�5/4&{��}1j�t��n^Ӽ���Z<0"էX�7a��d%�l�?J�*ǋ:oDC+���t��T�ƭY�~����~�_�U$��C�0g���
-���3'����L�OV��@ȸ�6�<U���Ʀ(�������h#j�w>�Xɓ� �6��ȡ�BJ��*�E�����p�q��R,)�5}���T(<�P�e˟�O�0Q*�zP˩��h�C�k5u�|U�����є�G|��&��zd�6����L��A��4��'�����I9��.!�?���{��6���i5F�p�Z���{��֩-���W[�@�V �}�ɐ>͸��>?DIي���/h�U�k�bUR��[�䗰�`�wU$�������,TǸ��R����n��)�)e]q{U����&��Tͽbcg��W�{�Sm�#�[)�t�D���[°��_���Ag�+�ɺ
Tt:��g���xj̕��b�}�Jn��{�ؚ�bu�m���ϊ�������ǻ�S-���}qɽ�:�nF�셣��(��f:T�*9����ٗ\z�L�,
�c���n������:���x�r�>.c;T\YB��-����rQ��߫�����R������(�-0�(�"�x�v�8�PI�ߔ;�"X��L�A���m����� 0 �	�s�W�b�*�N��a�+�}�1Ʀ$ә ۞pVi�Y��]ojAS���li4������������e\�>Xf�=��E�>a���k�B�?^f�knԯ�t`�}/��qc� �/0�ڣ�0�;����+l�}�!��4Ifzq�Gt�����D#�'��T�4�ͭ��f��5��YR�3X�fD69�⏔Ֆ-9�r�+e�*,�#X�?���01m��@7\C�g�j��)�ix+�w�����a �x��tU��E�j����޴u���Ð�#AB)��u�_e����`u��A�(t��m�k��>�F���:O���I�%���f�G�F>aal��R}�Qyǭl)�6s����]<9WaI�_g����Q�:)t�q��U��oE8y��0	�Sb�(ԛ�.Т�,T4L��4��Y`�͊�c
�[z?< ��?���Q_�������1���l�� ,�p��}ڏ�])v���S�i�(�%��Xw,+��օ6¿%�Ya	��NPb��7@������	Oj�GF�T#KgQ}TA
/)�4�z�����!:D ����F��(	��^^9E*�IU����ʐ�Ϫ���/Ķ��;���Z8V��?V�~L�!��3G��k�������C9g��psC���jk�@G�����;��B��ܣ b���t�3c�K�M.sa�0	?��l��8}��"�4�6��k{>sOAg�Y�χ�(�*Q�HO&昐3�B쎋uO�k���J{Y*rP#�f����Ҭ G�Ʋg��2/Rp�
����"�`Z��c�G�o&=��E��t�{�A`5+����sWEAFB�g�,��p\&��U��>?G�#��%L_߶����	LPZcU�N!�iՔ��G����@
��E���gq�ʚD��`)T�
�X 
4tQ٘{\�Sp��eSz���dW�� ��#M�RC��R�Ȧ�k;��hP��xvt�1{t@�Xw�v�q���Ql]-e$�ߞ<��sc������釱Y�ۣS���Fj�xga�OC_�D~T���E���z�g����.�c���0��q�*?��`��IT�X��q{�ھO��$ԟ��t�@#4ƚ�l#p0e�;��mi����m����M�W��o9��J�I���ܰ�OУ���SW4��G�F�9�F�={M8����<�5Y�)Z���s�1Ԝ)PO-��d	��XJc��V���]�%M�K�ˊ�>j����D%��D픶):Njf�ɞ�C;&�7�g1��	�%t3�s&�]](�Lj�LU�Qܿ~2�Ћv�X��l
��;4tĴ��B+7��lrn%{�I�?�lC�Ӄ�SaEnb�o��s�A��bDA?�]_� 'pHT���PTN��A�;�<�%�� ��@G��q�[S��0��,�C@��iL[>���P��nTLT&��><X�o�S����+0ܴ����mVh�l�����O����[=8�A&f`���3E�7�P����^P�K$J��}�i�����+��HS�	�, ��Ri,Uδ�"^
+�Q���0�~rqWM�
v�?f'~�4��o-��v,(�V,�ks�1'��=�-j���ꂼ<v���ib��~�=UB�.)�d25O����f�s"*��;����J�j�Q���rD"���!z�[]Gk���2�����(t�P�v�P6��%bn�%��Vs1	���j!�Z�_�շ���{5����c�̞�h��b.`u��U=�ir��F��1�z<:�X�t�m���ׇ���ƍ�����890@t#1��(��s��!df�?��Ϭ�����wF��� � Z���ʜ�_*�f��k�+����w�q��B�*�%hww��X��|Jw!�Zf�g�%�]���Ck�"|O��F�Y2ZXgr��%�t���4�&�����a{�\eJB��c�L]0��	���~It��������U�.�W�؆+���SOz��b8�����$5�g�Y=��������K$�>��1V=�����+:p#�JAY��c���9re�l�adhaw�J4�!o%m�ɦ�o�Oznx��Sޅ��.R�c-�A�A��y�V�Y��MW��ޥgH~&M+d���S�c�A�\q��}��,�R�7��<j ~�Lb����!��(26��4�<�~ᛢQ� /e9]Q�y�9V�{��9kO҄W�t�|#H��xy��]�PJ؉��r{ja5�Š�>�ΝJ@
����/�k8���UP;���Jnߺ�p����������sh���/�l�u�b�{T��h�5��g_��jօ��f-!�& �k6�z��-td.�����g� �=k|-@e
���g�֣����g[ͩ>0� ��f�Q�Ʈ_�㐸��b���B�	���7G:#��[�ݨF1�`�����%�H��v�fdކ���NI.�rݽ��I)B�'9��BI�>��Vp�^<$P���5jZ[��_`�{�?K��/౎�F+D����d n�9�.Ψ$�"$94���K�=_���vA_j���c�yr��Y��lD�3�6}��|>(��G�4l���A�j.!�.r��Dd����
�|-Ϯ��R��?��u�����
][*��"�PY��s
��4��랽.|zr�Qߓ�-ۏֿ�Bg��%{����ćX;��P�{�؜�ld��ޜ�����;(��(�\*`_�*�6�ϛ(�	�9k��C-R[�B�"ƭs�?�L�����o~R&9J�f���(Z�>���1$�66���ݭ�&X4p���N'h �hZ�
o`�=F�Nz'fă�0y;B`)[�J�%��NU^���"&��x�Q�����H�J�8�����O���7��q�썙��=��؏��d4_��H��uZ`i�����1��J�F�}ɄT�"I����i9:+`�����8LI��>q�B�i% | �2ˉ���T�MmI.a�φ�3}�F�bxd�b��aJ������]�����z;ɰ�B>�^\��i�JHc?����*�f�����;�ur�uL(;���l�Hǡ�����ʗD�� ���:�e�=W'R�y�RU:㨖���5�}'���֜!O��Oi Ty���kL�O�������ߞ�S�4u�j�����g	8D�|uFl�U�W�}jP�q�΢n+Gaqj���)�[�7U����O�!�7�M���ғ�e��z�/�Va*в�A�S��5����q�Y�� �?Y�=B��v-7��Sr�������s�o@:g5�2l0����(RS������n��u#o�j�<�NC����g�b�7]��bV�>7Wd��`��kH�4��#�;Ap9"�O~FPX�t�Pڅ�0[�}�5�1���[T���}�= ����!n�K\��۲WGE �8�ߡ��aӇ��=b��u
���d���ذl����ߏ��MH�q2y��ؑ �CM�f�0��u읅�ja,��T"�sR@����ug�y`��ڿW��Rۺp�gi>�il㷝�Gy��t��������;�lYCg�3w9Rg�qb3���M	}re�
��W��!�~�*���;<[c�7��h;�/"v���Y5'E$r����+4��?F��j�D{��Ļ�.&�8�o��&r�y�`c�ػۊn*
n ��BG�~�6�׳�%�("�5x�l�y��7ed��-;�T$�r,��oМ�,��lre�U��K�k�\�mB�˸���������4�H���w`eT��%����no�41n��0͟��7J���N��w"�5��PAia��]jm������)A?){y�h�P��-�1�^[9>�.A6u�i�=��%�zn�
|����=Y�,������n�4�#���L�O]=�3L��}6t�J$I�y!���v9}���ͣ��F�)�$��Ӻ�Vl�[�� \�#R \����N�2��\#��yU�� ��'�1��}X�嬯oT��tW;�WP�ɼ�[6�?�|�BDun�s庲u���,�-���=c-"lJT��!_�^R��I�׫�Q�'%���C�@��#�Y��a_�RjCq������ZZpw��6��f�y_�FáϗA_Y�mu��A[�3`0���7Tzy��d r�l.��@s��ӀʏF��mc��YE�ߩ��4�O��A�=���p�
�^�*��9��;w>e4a�����k��'�c��CӲ���C1q-�7h�^R�x
�EP�!ջ������?�����܏V,9�͈������wK�3n�$:�^�a3�Az���-0�i��'0ͮe�YY��I�m�����E�\Uhr�4%Z�a>�* �.�ayS�%�#�9��ê��	�H&���3̍ˠ5φ4�މV�i���d��U_���UP��V �M����m��� �ֈ.�ڊ�8 ��c�u�s��(�00�2����'�rVw(Ģ؊&p{M��=Vo����O�ÅlsƆ�����H(M���0�˲�Pntz}�O�N��]��H��NY�9�ŖP�~�Q�~e�C9�j1��C\W��j�0|Z�.�&^q���H������9��|�81V�2����mW��.�ȓ���T!t�0���ӻd`ɴ��v�u���w�(Y�ÔrV4 ��M�OB�����t?�CeT�H�\Y�R����Dt<�C�x:�A�	�,c�.�z��W�r��H%:��oy\FF.Q�!�	���yC�����U<��鼔���.�)�%�����.��*GF� ��	�Xw�
�r��\X�Q�z��>���XŜ�����`���-l2`�1R8�Y�v�@Ǽ�$�w��x�1��Fb){��� ݼ^H)��K��$+�9%�_��A���	�V���slHFс��Vf5R��{�Q��8�1?k΅P[�Ua��V={�;t�`���%��t���J]ϲb�2�*VH]L*e@+ �\�f�Ћ]]�{\��СQC��"��
鼧�a��ܔ_��3���/an�B���h�~�P4L��"��"C(2g��G_*�}�*�2gW̩�$��_@��2�]9�k*[�P��z��.����|�ݕ>�~���K��5�7�2����&~ 0�{6x�r5Q���8�r���=뒩����Osb�k:��c|���v	�.Տ�e�QLs��V�'$�p��y��h�]`�\�>D�ߺf��3{�"�s�aEׂ�j���3���|�hހ�C�h<�yҥّ�A�����>��	�T�N��V��s�Y`�P�g�!����}�j��ɵټW�za+6�(��8��*�x ��yC�#7��|p{�W�܍�`���=Dg��k����(=�ʎ��ip�f)��a=S���Ԛh����L��(P�B#��5���W����WM�u� �N��V_���/��N-���-�U6g�C��3~�^����<;��b��m�w��/��'&�k{�uf��$�ص�\�r�᜿}-�6!Bu3����4�uбv��M	�/hƒD�a�p�a"<p�'������u��HVپ'��0$�j��80Y�qF*�_��d�R��>�_jZX��7�%���v�CH����6�A�4\M����6�ܠj�B΍�&�9�����M����\�� ��G�aR�5���tkii!Û]�f�ㄿ��`ӂ��� ��{ϔ>5d�qF:��2Tw�-��c1��K^�<7z�
�Pn ǻp2ԡ�\v��ծ+C#�P�IQ�#,&وY���ɾ�D*��	U�A�Qˍ�ׁ�\5aA�E�Sw��]�#�o?��C �SMy��5)��Hj5��8p+�}Б�zS2�<Me�[s��P��:��I��sb���6q��]����ɺ?|xÏ��o�����'�l$o����F�g

Z��`g迕����F	}�s,Z�t��$��!
��:��S8���;v�'߄����y��U8F�@N��=1f�\Z,�&��@�c�ؽ�'��I�G�^W2�?��g��g�jռ@�}��`eQ�����n�p��s�Z���Oʋ��:J��F䀂lt�ʱ���=��#Ӣ+�/��'ndA��t�x8���xF8Ѓw�䀕Oo�	ѹEв˩�j�͂`�BB,�U�.�2�9��b0dbz�N��菚�em�����u@h�oK�{����r�)ywU�t9#�>fjdRH@~*�w�<�����a9$��@)̏(n�����ol���R�W��/L�B��/{ڔ�`_�]� U~�𵗜�kR>����l�RwHd�s�����������O�a�!e���`��'@x���T�f��i�&��|Č�rX�7BK�
��3ÿr�7�
t�fZ���hG��\�+�L��[~�P�DOg:�>�W�$L) z6��F�XmU� D������tU2��:a�"F=��'�㍱�j��h��
M�z""W�M3 c���4�f>��?�\e7��ٿE-ụ�p	)e�_H)�8h���%<�TyE�f��Cч�{3�\\n��j��6��_&k�����{Z
Y��#���h���`��I/�^�__��B��D@�Φ����g��.��3*%�_����I�W.��Z�#e
OV���ͧ��x�4�����k����)�[1���_*ހ�D��3<�=Y��	qzP������Xs_����	���	Ѷ�l�D�Nɍ-�8}�1wi����lG��$I��4o�I1�Y/�>�Grt��|ODT�G��֓w���D֗� _m���;'wq��V���Ad�_�qb�ݰ �{�n�k�s��t:�B�E,K�+�H<L��E��?����H��0�i�'���5���@sG��5n�>&����\�W��g/5�U�$V&Q]<U}�(��C�9Z���<�6l�����C��P�������6�_�>�U�y�k�W���8wE_i�W,
A"2�,]fm+�O����R�QhKa�S~�a��4�U����/{�97���G.��*J�aɨ�
w+�LH�Э#6��y<C1y0�.�W&4������㜈���E�Z����[>�li����q	�F����A>`��}ss9��8�2Ɍ(�$�K"���ddNrv�,߷�ȑ,&��,qo%��rf��s�n������lI�L8��ֵ�V��U�|��:���QJőK�����JgR�`E�Be9�oq���_.�\пYӡ�QZ�C�
�Ca|Z������\[j��꺷�ao���M�/��r�		���׃y]^ʂ��u#�f���m��D�[^�}��1t�]1��h��LA�;��K�q��mN^}�Y�.����c�W�\WMlډ�&�X�mn�G%��E;>�w;sj�G<a�x��w'��c1j�����u2�H�0KQCe�@�R����Q/)g�C���-b 'z#��Y�P��ſ��U�P# �y�k��(rG:�C����+�>$�H���u����1[k!����h����ީ�z�	�W�$��渃���0N��M���^��VNv>k�,F��Ԙ����إ40�I��k��Y�g���ߴޖ��1����I���ЗP#$��4g<&����^����*4$��#m5��b��$$��8����w:�u�sMGo�~��������G���)�s�]��GV�z�L*ކy�HS�_���LK�@�=�j��	*uڣ�_O�����T��H�?�͂�t"��Ye(Xq&���(�T4)��xɺgy�9,��%͠�t���/"(�:�=�owc���Ckl�[����/�����0�'�A�?�6;##IʡI���� \�h�GC��_����4.I7���r{�SX��eH\�Q��=�zb���8Q�x�$P�,*b��}��l*�ǜ@xLK3���ح_�����2���@�p3�OrQ��cd$D���Ypq�z�����C7�H�5����KEӔ��"P+���AR�H}��}G���'�>��t��x����S��2������_
�b��J�+	9L��tBB-(���2�":Uj�Vc^6i����8Jm/���^�n�6�( ��63%�C��cI�5sJn��N�� �@�ntc�D�&��|���<�E<!�0d�(⩖j�yy���;e�qC�vP�7����(~��j��_z���T�x����d7�6�)RD�"������g���E�~ ��ȓ���#�*�-a�Bۘ~b����̦�V��"����Y1I��|���^Yd���-�Ye��Ȳ�^���z��������a�ǡ4�`�QX��_�9��&�p�����pt�f:�v�f�A�c�9ʬ�R9��5=x	[G�R�6���8M�G;J�}iB.�B�l�	�܋�	�:ȩ�@��Q�2���!`PSC�?��;�6fo����聸!�uu������4�1Wycp+uW�8���_}1w�?������F��������pq������̣��_����pL�e\�y�Z������L�W�Z���)�i!�X����A�^����m B�]#��׹ed�`��+�F��m�2�[�)�7e1yԲ]G�!�sX8��3H,�w��ż�%.�����ꡁ�K�x������>4Y��\"��8�F�,4J�[nV�O}�Ktw�>eK}u��B+5{�7�������1�	���<�W��,Q�����S������5����V���?�����*vs7|�+=q�k��/y�"ǅS��l�A�U&�7���	/NT}����Q
�s�c�ە�S��	#���8 �����t��;k����Cb�����ń&�1�  � G�$$�t�pt��y���x��4)o���c�;��M�9t�;6;�sC����R�Q�|I�N�gNc�Ee.H`�-7�9ڙ�x�-jK^	�)ȸ�qdH�tj��2-��i9��M�R]�ԝٟF�g� ?p�	�����M��yiW�Fz����J�E83���(a�e�ݗ�����������;��M��P{,d��.�<a=�{�r��]�@p�.�����H��{�0�A}^�c�f\LOox\��i�a@$��"�(��J�
\�nF����x~���<Z�w���)��aŵ��2BL<���X�mxIeU���p�\�\�O6_�m]Z7�+=��){���1�_)�V�� [$� o_�iVq �w}k�ޜ�����55&8�3�|�h�������$�^6�P��SگT���,�hq�� �Ũ�&s���mЄ#�kU���B��n�n��������^l�ˈ��4�Ρҿ\��r��Mn+�~{L�m�c�SJ�Kߧ���P���|X�Ќ���hR�u����iS�;Ó���X���D8�� {�R?T����	HsW���]�>�ky�o=�+�[�[��kwp��B�@��E��Ƅ\���*�9�F<l���Rt�1#�N���50jd�[n�-El	\k$��5Q�8ն1HF��J���p4^���a�L���t�7�FkQ'c�jgbwYU���[.����U���Q���ft�o�u ^Fy�V�O0��
ZZbB���7�*�mQ?�S ��]�ye3�_��@��}����F Ͻ�ȓ�@(%3���kq�}�	xo���Qʩu��2��~�^�\}��hqI6�H�.)ɣ�r���[���HY�)�P:d/�|p�����$,�>	C� �<K�����N��1TH@g,��&��闠9&��Ӣ�ꄦϵQ֓X(/��K����$�o�w~b�wɿr��A��Q�k`,o{�  �_l�����Q�5�pw��"K��Rhg"��0���.�<�Ӓ ������>�?q��"�*�-�т�B~�X�m3t��o�8�1yY�z�����4.?c#�{-ø�m|~����ŞNI�m�>�0
 �=�G��}�$N[�ճ��.W��k�C�(p�MB4�T�D���xe��k��ͮ��7��d��a�7�|U��wl�f����r��81gUX�ԝ��8fKT{p�̟*���U�j�T�e�r���Ib�Ԃ�o2�	�p?�$.�O¥]Ѵ���C�)�2����r�Ÿ*:�H��d���.*�y�����j��u������z�HA��']f��e�@A��K�h�m����7�`m��L����������_���i��`��A��}�>\K�j�*�Kv�%|�3"?�gnR3�+D�<��o�1��p{o��t�\�H�䛸����lG�&G��^�B��N���
���&�%|I�GYy�.P�ݰ��>R����hY�Z;����9C7ְ#�'Hg7.Q�3��Z���5}'c�"��ZQ����!E�:��+��J��܏d���y�He�`���3�f�c��v�6�;�עAFh	��ta@��;��.�*h�e�myv������R�"c����S����ډ�.1�]	|Z�&�׹�wx�ߎzKB�[.~2R�����L���2���L�<���v�-gE��$��w�A%���8�0��q���0o)��"B']�3�ZY"wDT��������*͂�Qv,���~�D@`D��?�������$�ږ��@^�{zu�I{m�h�;�����e�[�(��N���ۂҦ�<]�ʜ`)R�ͼV<td7b����%��eYs�H�@�K��hr��ɥ�$��#t��-�#�X���a�&P�N�ǎ%��V�'��ߨ��9tp�["sʎjdl1��7��l/}�A�*.�;oN���}-%4�=wÂ��[��}�7�h��V�j���~��VՋD�%�V�� �{����c�����^^���ü]��7�Zly_ҩ9s9�UV�Mch��*�@��b�"���ҥ�#�6��h�e���e򚕲u�na�`�֠y3Ĺ�yh.�D<߷:z��*"����d�ѫs ��s�I�a��V�p/3%C�`R�ؑ(�����m�̑|�����%=4Ͳ�Nh�DX�'���5\�a'+������b��<恠��Q#�>���
�u?
j%�n�Q.���8�M�e���1�)H�w��~Ey�c�4������ne�&oxi��Y�3FY��ه[W$;����(�P�C$�^���dfTe`����Lҁ<}���ENh��d|���=9_�'Ɗt�L?��(��wI�aw�u4����rM"f3/��S�5�l\=Q}v��5Enz�p}�ੴ�Y6�0�V��z�@��㈝��S�S�=���Q[;?�F�bg0%�U�?0s�{"�Q�_Ϳo�^H��_q'�_�	ZF:���b|�|�{!��Mu@k ܫy���/�p����D ʔ��<�����(��y�A�{�fE���(]�j����޾o��2�3��殺S��Z�P�" $�S�\����4�~���Mו�삣�]@����}n�vQ������~�7��1�.��	!�#&B��C;�eD?	���]$�1����	��|���޽=念�F�d$+���0o˕ڏ&4h�ՠ7,����˂�Ӈ���&�_R�wQ03R{>0�߹�6z�D{#�hn�_-A]q/�_=����x$�@1�Dz�R�)Dh��6t�y$ ������!�Ixրk?��-8*�lR�;�!c����^U���NL]����.�j~7�"�iMk�T��C%bJ1���J�n�e)~[�
�ז��!Z1t��kHR��Heu�ޜȯ0���8����{��ВR_>��HԹ�3�a x��K��E^���~)5#���4�8t�g�,�zN��ȏ8.1P,-����ZSLr�~um�?���7v�h<`������5��4��u�n��}Ʈ�w]k��B�l	�������=HϪڮة��W��T�?c�G^0MI\�C:`^M萂 �5��&�1�%�2glz�R���:���TQ9��(P�LV��Y�1��j>���E��{R�G03*�fT�jPy\������Q4� ����ie����E�}������X��d��^N���t��'c�?��c��hz]�^����U�Z�'��c�<y�Ǟl�4oᷥ�J$;����z���fxi�X��Y���J䅣q|�Z���m+�`�KˬN�%aõ��F�Ò_�3����,�"A�Y琶$�.�L~=�yXQ;#��#�O���y��g��*�.h�����5r�Ą�3�'�4������ƅ|��_.o8/*�nc�Vg�a8���	߳`��{��!�̟�Q�BU��U��Kk�2' ���B�^����!?��W��Å�������Mس��{�b�����S X:6~�]��[����V�j7���Mί*w% ���t �d���3�����<	%Β�1,�����"]O�p������������G(_z�Y^�(��q���<�Ƞ����R��̰fl�¨���ƣ��m�6<p}[^z�p��;�l��P�]��a�?U����\t�X1��w��_R@���93��E��{�b��b�L��/i�њ�@�D�����]`ɾ���I%�7�.+Z�$�����f��;���$�*��Zt��-WL�k�:�MG[G��t�0. 	�I�5O度�'��c���zm1I�����FϴlX����x
C�Vل8�A�	��4X
:t�����0��+��{��7u�੍��M�nz/'���3��T�N)d�+�𵋷�sP��(������7�iϪ<4�����z��d���N_�v����b'Q�+����`����u}Q��B�o�i�0�����ؠ�}�dᔒb��������G�l)���-	=rɯy0�]�+p	�����PA�"�UЊ���&���r����~T���H������m`e�N+�uvn�����#�٩I	4G����w��4�Md
���;�G�icXs�\Hc"@#�����,�� BSj"Waak֙*i�QD��p����h��9�v=��8f5�`Y��^���
���M3�t�J�Tj���D�w~O-D6l�I����G���m��7�{]aw/*�f�ݦ��$X2�eWU���g0����6eyj���У�uY^F��d�\;�\\��kwWRk�GHAQZ�>0VzbJ�g����8��Z� �ȓi�����O�~=��h� ��A���@o���F��M��T���W&xc�y+_��8ĥ3����0��O�C$y"#����m��Sr��[}c��-�,�ݎ^��P����q���z�\�LB���d�\#����u�Ƹ3�e9Sq�%�B�K��`�" �Z��= tL0�<w+��T[,�B�vj��*P�7ٲ�9��Z�����0 "kgx^=B�Ud2D��t���I���I�W�U���ܯ��z�:`�f[�����O~}�̠'��e)}�f�������Q��(���r�}���_0b�Z�2���# �9�����J�|-�9�wBH�z����Dl&�	�u�=V��9� x����G0������ɢ�[}O�M �^��B�<�?�0s���S��Aͼf�q[���#Q�4���Ν�0��S��F�F�`?-�b鑖F[^��*vJ�	�ױ{�����p)Tf�o�u���pBP"uE�2�$é�Q��۟^�]I8�^�|��H�����;8L�_�\�� *���7�wE#�ڜ��������!�d|���_?,W>1�E�]ym����m�\d����n�e�oLU��o��ν�=>SX{[Џ�cz�;���D��9b��)�7Q�Ǔ�J��\a�5�����g��:�u�m����m:�b���p��s�z�tL��XJIfلP��CdnBҴ��Җ��}k����M��K�@5���辌���~���b�i�s�3�pk���daj��W���i@kA�1}���,(؊����� �����R����������� B���֏��O�S�2��W��z�2�%��(��'����3�w����$�C�d���"�K�MV,T]�ʟը�=x°@�b^��f/n[����5Vo3�4�M�����]]��N���N��Y�y�0�dl'0���ӎ|پ��D_Y�	i�`�6F�.\R#shI��t��h����NMӚ�|�b�<��B7�H--�2�,-�v�N�Y��}���ĥ���G���b����I< ���5����ߨ�b�o�9��Gɩm�m�@;/ �kn/9P��Aصz��11r����|oq�RG��`��#}�gO����� n��h��_g�\��|%�KЗ���dX�]#�kx�6�J��$���mJ�4��|�O��C�
:b*b6)��0C�်	3�_} �|b:����_H[�>z�Oh�薭Kt6�sk�U�5G��!z���fDKw�֨�9s��`V�*3�f�C������`(��*��Q��r/���8ʧwO�%�+gʼ��P��|^{ ����&xd�qo���%���~l����	�l;�L�տ��Pr�b�)L@|��]�b�ߣr0EK��;�kN��Y{����j���.Q�!��!$���)9"�o�Es�2@W���d��L����M��+��x-W٭:D�E�@�U8�� �f_$�v�t��<�F�IT�mE$`U6\>->��h�y"�#�BDѴ����P.S� |�j�c[6V�J	�JP@�d뢇��C`~�4������i��R�#,7r�~h�p��-��Z�W�C��[R�Ǉ���s�'u1��������Ӑ�� ��.��b<��O�h��<O�	?{k���Ĥ2�"�� �
��ܪ=��:{�|G���i�!���¢vZ)u벃��F΄��� FZ�W�vb�a�Jv���=��u���|i;{#Vȇ�Y͂Y�!�VS�/M�hUn�'-�O?���;���lJ4q���������-�kz�� 4��Xz�n`Vk��
TZ\?!��}>�3`~���i�P@���Y�����E�ꔿ�pO���V�nr�s�j��{v�pSp�=�s����F���BG�C�V�^x6Z�� ���)�͸a�A.Aȸ(g�+���X"l�K��o��lV`M3ܕbݲ	�gT[.�Yp��0U�xr�	&& ���k���%����,�$�S�,T#�Gl��2����XJ�?ߞ(#��A����ꁝy��p������7G�qBGX~
���7������2��|$�iZ�J�6k���Ψ
�=X؍y�ż��ԒN�?+���2�Dk~"�&��b�$R�E�Ɋ'��@����5I�tw^�c�Ɨ���E�wQq���R��w���΋����O���"O�a2J�scٿ���װ���XqD��K�K����غ=^�b�ZЃ�Ti�]=�d�P�L?�U8��G��p�Sd��">��p�Y3��!���;�غI����HZ7�l���:/�*���f���N'�	���o=��b�C��	녕ᣁ�����[^(���?����� h�,�U�������}~8�i,,�ނ͜����*�m�x!w[5����K��gO�IYDj�C�C����٭��>�K���?JáV&����1X���o=vev����⿵�	@w �)}U{5��m*�P�+�Y�s��o%a�U���ї��6�o�ILy[~��%�7D�vA$*U�/��.8���($���)�huQ4hƓ�m/�[g�,�u44ES�Pې#�b�fs*��B�@�MG~��>hh���C�a��
��a���uB,��G�Z��s�!G��ҹ�3G;�浪1p<~�� i��
I������`�J����N<gRf^��6s��[�J�%Jw0ט�]~mkz�A|���m��&Z�%k�wF�A��u$=D+�A��Wxv�q^���s.ف�9<Z4B�L�|Ry�q����^�Q�����渢d����7ꆆt��>fV*��N���鎞퀋����E�/�<ݍ��Mog�8w1�Y� [c	8�G�nz��s"��Σh.���%u3l{lUQR@�����/\�A�6�N�'��y�޷A�� �'|ږ7�����8�4��=*�~�Ձ��/���Vu��ώ_Yj(sk��< �,p���m$=��WL1�f��� $���n���~��Z�
3���Te�ok�Vp�]��XjT��S�z�U��J����C��s�� �h����K�m\�q�~T�,]v��~Y�?8#9H��6�X2Y���3�3�)V)Rɶ��.���h �i櫭"��.9�[Y�dA���o���T�������9���ǒ=;e��e�»<��@PQ>��jNV���Q�o=9KD�)�'Mõ����{�	�U<�ẍ�|w^k�e��%Pv�g^�Y"i�Y��Hî%o<o��P-v~;�Oɹ��1zl@��E/�iٲ�AfP���I�?��
�6c�aJ���u��>��t�h^�ߙ�2�p�(�R���"��]���F����.Iv�����ԂE�ǰ�N5��6�	 UB^&�%`-sP��l5A���f��M`�V嫿��ߔ��@��h�����\�P�	�!�?����ᲆ*�ڪ������2)7�]9�B5����a>��Y� u��B�$�hl�����t��}�7�DO=��f�3qz`�enuO�S���^��;5[)��}�4��ğ4�{n����p�t�K�-^�@|�9a5eS; ��R�7��=� o�8��X���7�}�����K��dzm���Wf:n�l<U���Z�F����9ܧ�!��0N��%/��:���� �0�Z��s�����9�,�'���[�r�B�9n>��c��(�4�)�ͽB���;s�v�����i�}�X_�_��.�Po�׃��`z���T��ZJn���za�c|�e��>�٩7��m�tݞ����tA5E�`P~����b�Fl	Z�����ăհ��>�L^��B9�j�z'?��@�(�zD_�>AX�}9�v�x����ɓgw�^�J	-��	:Q��4W+�O�BP�}b�V@��('ߢ{���t3�.��@bءbyZ8�t��wuKl0w��2a��B���<(x�'}C'����L-t~NC�H���% �B֗E(�;���f��#�=�?#4B�1��$��6�k���$�cZ��Kά2�dP�}�"E��	����K�2�%���"~�e�/x���ߛ+�
��f!X>���&��7�+� KJ����uQ�|�����T=�5?!4lF?�������`j�l�,��㪁U�c�\@_~���[��S��Tݑ� =v���h(}\|E�%��+]�;��G�%�+z�g��pR�k�Xe �=��R�N(W%<�ʌ?���pf��P���oBU&�gG��?1	Z��ꤡ�ݙ$��$2�m�Q�r����exR}�1z��~0lṖsq��߳I��z������*(���,9�|��*��3���.ZQ��M��ܪ�GA����_M�C�Q_{fՄ��կ�|�I�݃���p�#k���,�ea�[��f��s�$��j�쬀
V'���K6���u��G�>Y�ר ��i���wl(�M��+�U{\��Z`�e,��:�
�Ԇ�
#���Zi�L��Sk���h��I�0R�-ڨܙc��/�	����A����bZ-�A�,?!����fnBM`�t��������-�h�0rz/޼tU�w(N���O�e�����5�W;�ј�k��|Z?`|���l���ݗ'�\�@כ�c9�X��fW��S#5`��W��w ҃s���?.f}W	��`>��O?Hc�0��[�DG,0�/�.�|.V+h8�X�h��w=!Q�H��vp3t��V��0E�%��C�3\��d��&f��������O�۶�k�g�V����/���ssc0/i5s��#	��F1���]~���:)3�4S�U+Fg[�/$Y�	���`�4y"2�G.U���2� \�����Q��j9|��<���y��H]D�!d��M_����֏_�4̿~
:��~� e�+�u露;1Ά�"Ca��i��R��l?��Or�R��\����Y�
؛q��%˴V�F!⡸!_Ľ��Ł|1��U�00<�ԉ/��Jy�VIXG-4Mk��+���V���8�Ƃ���nGs�k~�q��-R�*��O�-�"Y�;Ԛ��c*�k8!���[s
��2�{�oUP��e�$�?f 7�����kn�8�R�/\�֏0�U�����T�i�7����}��t!�D7����2P�DdJ�d�IfX�i2wƼ�4W4�Z��]+��٫I��:�nǂV���:�&x�R��c�S~��Q�9䩝���׵��+��!��Q60π����A�[�?7�RO-YE��ߗt4�Z���֔�j_iU��#}R��ܮ̈eGa>>-�����E�">֟�n3B>�r�#gƪCl.D�A�d�^Y����9E���Ϋ��C�^xG�S(��$�\c�y���YWyX���ц@L��ـ�[�k�d�hd�f�/�.A�@�s��g�4%{�z�CNGIP4=��E��<�l��߮T6��Z��fa�d�U�L��p�t�qR��n�҄U>P*�pI#9�٩��c��z���}bt�*J,.���~��$��Q}a�JE��?-HFQ��y[�;����:����*�<�L�@�����*#�>��εm|�JT�4��a��[z���VS0���ۭC�ᑰ�?!�O���<�凷d	���z���<�^��o"���A�.�T�
Nw1`χ	�ڗ��Gj��H]v���DVhޘ���e�&���oD�zW��&6�q���@5|�%��gz�L|f��8!@D�%F���L +��`]3u���˒j��L��R=X+���Ix�S![l=��V ��7v 0Fc���c'��_�!m&P��mi^�)%
�)@�o���m��l�֘]�dc����E7�w��n�+��3��)�݁0r��Y�� ����\�U��u��j�(8[k;�&J�X������G@m�Ѯ蝭/�&%�ߛ�1��8D��ri��\q��U]#��`|��s�m(��;�F)�<rn��E��Xxt�WjaS���G��$㷚.ܛ����ʙ��m]���P�{y{<�!�D8 ¼�x���\R(�k���] ����p�6��_������ �Fm�j��}�<�Y��.�_�:X@�e5�rC�!�:��شo ��=��;b�������u;y|��@B�H�o��Z{�:�/��Zܪ6+�M}���Q��9��}���U�o�/äR��	r���yI�$ROWv�}��Dp�No���#K��?,���������$s3��9������D�豒��i*��
�x\ɶb6yW˞`�4���jS��ky_Z�3x�,�t�w��]��z��~����఑��`�oR_�Q�xͷ�	�i���35��1�;�@�9x�¶_����ϪJ�O�����X�n�'.�~Z\'In��Z1��LNn�W�p�ն_^;C���`��3=�8M�[�ܖ��I��z,�!i)l��C���=i��&쳏��[�[�[vn��wdQ�nރ^��(�I�r�Z�R��s����4�Qq���,[�E�����ˀ��	B���������j����p �v��^�ƳL���4S�a�\sT��qK�[(�F�3`1��\!n�����}��(��(�!"6X~"�n4���=:?\QTG�*�gr���/F	Kf'��	��T����ƪPE;��\��pB��
��G����\	�����9�lr���^bcR@i[�7N��1��Fzfe��P|7u�_�c�?������R�y�~�ׄ�fw����{�ϯ-D�̉�3�+?�PtT�T���*#-���O��up�w�P`	wF7+S��|K��}ԟ����j�_k8��V�Th���k5��B�4�6F��R8TE	Ec�6p���T��x7e�Y������g���1���6zKq/��C�]��5���UT*��F�%����hL/._��ei*��~G�f�����2��;�dr�o�WZ��S��ć��f�`j���;ƈc�3W��4����?��1��u���M;�o
c�y��H����6mgf��T����=e����H��d�F�5���c�W-2ɇ��<
�r�p��}��N���1�ۆ�T>}ٚ�b��6�~:J�^�V�";��:�������T�{]����*q���퐾�zZ1�$*�"��0�F�"ZZU�v|}a�$�I��H���Ly�R;��� �����Ush]��"�XY%��5FE?�"K=�j`�:×M"\�6D(��AQ����D�(��2S�H�(�{	��N��3��񶕷�����JI�E�=0S��d�]K0��)7e�%	�0��-W��1 1x*��;��7ɫ�l��R��.�{1�4	��U����e��
Θ��$�{�V�$0�����vM&�B�R_C�x��!�_�"7�H���&]�:D�B�TT��B��V������+ux���YէO
$,s�:r�.@-�ه�&��F7������(2Տ��7��{_<�J�U�������檢�������2�#t����G> 2��eѮh��Yʫ��Ȍ���XJ�\1G �_�^��� גM�to�7u
�E�q~?���
���,fTW����4���B����G[pDB�+��ҝ�
;s&�[^�l��*O��=<��GS*K��ό�e��#I�C���f��VL�9��gi���$:$J>�<��P{TF�����-�ka�w�ئ�ځ� kK�G��������^��o����y�E�p��ƭVM���-\y^�!39�~w�V
�*��G���g%iY�A1Or�JF��i������F�>}�nAw"y�}��Sq�-P�%�y
�l���K��i�I���D���ʶ����5ןp ��I�1�H���&+�5H�g$P��{Z����p�ӜW%��f�ȕ�k6�����by�S�QM��H�\�F4{���1�=*!֘�M��з\jR��5c�+�b|1�|��R������S��|Q[�"�7�f�""��uu�4_Ԭ������sM�1L��ƌZ��X�L��m��u�'X�aj}�3�k��Z	��w��a���8
��t���2JC��f#�;s���{����v�wo솔$��!���*+�V�|�$���|\�C֟��(���)9�W��ꃄ`'BօߟS5s�x�N&�t�T�c|q샥��E����"���y�?HQ"�a�+�	�:�VE:ʸ[��� ��u���7O���(i,�"75����W����u͢D,:0^���({ 8ݎi(�����՛���X
��>X�,c���	�~���k�ρ~GD#�׋z��˯}-�1�)#(�x�~��B����/�s�ʺs� wa3�,���lh'��nP<O���!@�K�Z�G�HU� ���tP�G-Ĕ ��Ȧ�+]zԞq������]���뺙d�ؕ���8M�w�:f�y���+��Ay;C?$�Q�F��P=[�^ ��[/��#�Q&,�o_���f�b�r	9ey���.@�Oe��!��!e�E~��"�YF�L�����C/����1���9�Ӆ���jY��JO��?���Y@^�cEٲ5�5�!�_�#�9��d�#����^߹F�@E#�ɯ��#p:�2�9Ba�a�u4��:Z=M�kՙ���=#�u٪)ǭ���@8*o?�f��3s
�?�Q���F�t �Ƈ#̀MPFǘ↤�ۜ�ek�Ty��>1�q�/�-� �m��y 1��i,�[z�,�%�j�Ǳ1�&cE�7�j �Z����ۋb�����lh��_$�-g�F��Q5�Y;W��."x��`x/4��DXnr�;��!v?%=ذӄ�gb�Wv�l���E@� ��~����in[S(۬�H��(X��|^�튜���"���m�~�$��.�R,9N2c�J6K��]N�JL��v4���S�؁e�Mo62H�]�S�_�yD=2�\@fE�r�D �'e2.�<�u��,s��ɲP�RBq �&.<�����H�I��x��oe�\���4�E0���N����D���?s��5$��I��%��7u��w�u(�$�5Y�p�hW)ya�;Ѳ�����|��P.���?���uR�cpܬ��GO�o-Tʧ���E7��'.u�۪o��n�C�:�Gd�j�t�YH���J��<0�{G�];��j)d��☷^��-ޡVB	3i��HM������\�XZ)?����/9a���,RE��ӗ�M��Fs6��4jZQ]�W?� ���=�������1$$&��^�}�a��Vu�^�L�|�CΠ��!i|w.-�]!tɀA�c�!���4���\�����X���'���B�<�'	��_ڴ�賎�=՚|��ҞZx!Q�c���V�����pq*���*��)��,7����q��"@6*��v�$}rHL�Y��-�ɷ��Tv+�u
0�����f��gUY��r�1n���0G��9vϭ��,�4tdn�%�>p���*|�27�]�֥g���+M���Ō�y5+��5��p�����!f����hm� u�(�N��b����(e.�p-�c xA�C]PN�� �N��+T�S�o0%�Nf�BI�K(A�yҧl���cZ��FDi�i���䤽X�ך�
qT���!�Eg��\�H-���H'�ˌc����9w��#T*��#�Z�R����ʂ������{	Fw!�{��#�F��*z���m��N�WyQf{�Y��S�h@8�К����\�up��z665�8L�U͍�r��ɖc�	�%���,Щ�1Xb��*�󗪉@�(��&���шRCyN�"j�.��cL��c��i��4��c�Zu�q&��2b����H�*�[�E���h�lCu�Ϡ-=����1)C���L��rsϓ�]��H����!iIu@���L���o��\vP��(PC4�j��{X�gVt#�F�]2Mb�^=��8��ޫi-�ټe̤���E����L؆��i�PG�w��p��F�a��LzN$ڥ����vS����`^�c��k���C����Ă�)�A�(�6@��[�m#��F1���"�L�d<��Ϟ�͘��B��)]��Y{�V#��k��-F)��ĕ�F�,��\�G�pv^�~$���1I�=���4c6�P�/)>B�)��d�r��d�R�O�dkE���,{q�{�J����w;��k�vQP�~�,����'A3���o�/u�ߴ�5��c�ut�*�2ttl\t���6��>^�K�O;H��z��ѣZ�Re�� ���a7�)Y���8)o`J^�����,HS]c	��9�z�y�hy.�����ݧ���^�[f4��?�6ޜ�.Ѷ�v�8�yi�P/�wuH��l�
�5>�]N�mrL����Q���o���@/�v��M=�"/a���$(�W�V8��m�٢�y�H��=`�JJ5�[F�ݵ�ӛ�+�@ի�Xu2�#s�	�Q����#�AQ0<��yE�~S�q<kh���'��Sz��ϗ�4�]��k��Kc� �1�N+��8�TV��4��jg�Yz�գ�Ë�*3E��a|����y�f�9u�TpTܦX1��T�P�bi[�����Y�cԲҖUD��f�٭=�ª�RnzT�w\�?�E���Ag�ϧ�FZ�J��沇�i1(�1�V�P��}喹1 i��eh'-��X<`N,"��uדas�����J�1�_c7��<���H�s�z�P��蠄m<;W��'�=M�>!+@�I��EMVvf��no<w 
߯7�x�rۨz�FhyQz�}f�-����6wx���Z��������N�[����~DR�cb��6{(=b�2�比7�S~�T��F�$�c�(�a�ȿL�!f6�Xk������u�rSI�R���B;{����v�'�	�+�h~;2�?/9Ø�bq�7�Rɚ�|D�A
�B|��y�_��e��u�;os}�'�!e�(�Q5I�XAu��0.��=y8N�����J}��)#���&�b�b���Q��<s	=����d�{��������H�ŉ:�ԶW8�i�-�Fv��}�}�s�m��E,*�B<y�GMIj�H��p���v�����"�Q,<�����M�0gD��{r;0᝸`�z~q���2��O���$�����Gy��	�O{�8|�SNOZ{~�M����	��,������ޙ�M�-��>�$IJMZ��__(�MF�xNIb̧��ኔ�5H/|���m'�{�_CAoRQ�蘿��hxI�s�w��K�K|��,>�1�1���ͬ�Z���7G&��~�9��e_U?xlN�3�-�KĖ�n*�%BCIpX���-:X*ibva$Q
0��D���]̚���9��(Ƃ�0���K�?-�6z$N9�o_� ���n���t��je$�r�m����O#��@CO��.���R�����p�ÛW\N�'$�b�E�jo�t�l���iaA�}E��6���K&:!�$h�+��L~ز6O[X��-�Q(��BQf�Yv�/S�q�v��U䢠)e��]�	ê���S4bpN���~�20-������ыF,��9Qݣ���KN�-��̮VH�h(՚,��̆5�L�ْ�4�}VM���HY����(s ����b��3HԥB�S�!nv��u�H�ߪ�r��}��7�S�lO%�nkrg�Y4
k�}(K$;�kK/2a��=��̾`6ˣ� c6�U��'$�jClԸ ��6��P���|5,g��8B�c�Q�Y|9d�%�s��FrHӷ@*�	�U��r'|��)��Wԛ2��C�& :GajTte�7��RuG����.�^:��rG5.D�W���^���C���gT:���w@�����7"(�
�D�Ir���CP���th�|�ƣ�\iqY�����̡����������D�x+���oW-O
�ֈ�6/�)�2ID�$�%��+�I\Mx���69J><�j�J�etO��?��1�i2'�s��$�L�2ڶ��f18�l�"(���]���	:��A��2�:�� MI\�n~Ս��=�C�F�z%:s Y\�Ԣ�,��w���Xr�[�� �)��M%��)6_��`��>�:���sa,ԇH<̝�	�3ه�,�'����3���`���h�!˷m]^�l)6� 0vb���M�~ؑ%#�^3c#�����c�	�?����ʈXf��O��k^j\L�H�	D0���u_E5Q�h��61�pcD�-~�i��㙍�+e!��#�	�	�2��ؓ���&�A�c���~z���E�N	yʜ�Vɱ��JLb�!��uUn�t���#ª[����q�����0|�9�$�t����p���C`�����Tvߙ[jH�ɠ=lg��;:c�ȸ�&f�к�	����j^���E�و�N^>`c���c����{Mn$���5�0�:�P5lii�I*���
)���5���{Q�2��`;4���0!^W*uҘvW�<�6��~�˱6��I�%�_�8�&�j?ơ�� ���{(�[G�8�0�C��Z�N�����
x8-��:�'s��K�!Qa�����5��Z�U��y�Lr�W��?����W���l�R���18�^ˢ���y�����,_S����ݡ&lR�O��j=7�ۊ�\����S�
*F��0~��٪^#[�et��u�/���X}�o�X,�B�6�T�}A���+��U$��zc�[o��.��P �J���W.��
������%��Z*f"в����|�iF0�H�n�@�Y��pjύ����+�����0�2�(�D���^��Z����&@�f����}�)��2\ĭ�I�{�}�y3���H ���Ay΀��g�W�3�-�#�>�G*�߾pB�>W$蠹�ڕ
9�ҷ�Y�t�D6�+l꧐�Nh*Q�M�0�����iM�z���F��}K�Pb�]���&r�L.�>���b�U��t�H0�f��П�,3�Ց¤��3&�g����V
PY�`���7_��S^��{�W��fnE�5�*�5��}L;p;�ucB0<�Lyq�Մ>h�*T��e�{�%MϜp/��@�/��`%�x� ��g��n�&�ȥx&���CY��#(x�4 �ɕ+x��S  @���{��O?��ƀ�|Kf{_�(�"��FQj�d�ɝ��D<oH�!����7�F\|A�3��tGd_�,7��1<R@�!�{Mt*�������5��6��GŎ#>�mj�Y߅%V8��>��oτE�_��cG<f�7y�Px�b�;JB� �Ŝ��Y8�H�Lg�|�.rw#�ͭ���e5��8��:�_�'%-&��,s�/�!�3�N���-���ܤ>"��8Xؑ�-��w�/Df}�
�~)4|���)��[�n;0-;�&��T5s���X�&H���Y�jW��'���lh'��X؂���9�-����q:�Ⱦ���S�f�5�Q,�G"eN��]=j?5��؟�,(-���Ԏ9�x�O��#M;tp|EF��t�\����|���n��͠��h�|Vh�*�0d�;s��l��Mz�5|��|�𭏿�7<�����G
�c'�=^�N��ht� ?V���Ƭ���2���^��Hg����'���!�����3����Я�+��oj�K��V߳�T��R�0U"^ɾY2%T��F�|����Ґ���t4w��)*�[N`��g�[�c�Ad��Fhw ��~� ��|�M�A.�x&?��5`4�/UEo�FWM��!��כ9��[xt��.�/ҳ�%+�����r*�jl:�>Cs���*��%�w�6�vRo�Ry�3�`����?�1��j/���H�l��5A+�u>�h%q����F�j�+��BV���N�q�G�9�ʶ���*�-���߃x��l9D��\F4���7xͽ�e�Ɖ�Ed�_��0�>�i�ԭ�$�?��1+B��TYP?f+I�D7���ʇ*�o8���I��'����T�:��)�T�B�Z�]X��g/�J�X~�겍����B5��s=d�8YB�Gt�ۣ���8t [�@�)���Hz���ij*���.���ēIQyd�֯v�i6wF#�~,�w������L\�
���qCL_a[���t�+P7�C�Տ�������f�x��O
r�!�W:YQMh�3m��YΆrrFI��/�r�s�P����B8�s�F�vϓ�t7	ȟLt�1���� f'a��fd���:�?&��Dݓ�RL�[+eR����*�'v�?:�/��zw��|��j���Ǎ���A�S��rt}��q��~��ky��Tm�h�BJ�*W�=�B��N'*#j��E�SO"u��m�2����@�[ǻe*�rK�,Ey�8� 88AJ5����Uf�&����l�����S�e�S=`�_q)��_=�hq�+�{��h�y��ȿ�f� Hu����B�)⍖���X�7?cp�$;R��&ѧ� C��m���ɥ��j@甕�Ʃ�¨����/<��P�r�w�`zެ�υ��R-���C���	�Mi��#кx��mo?B�x��䰀�<;�w<������4 34 Q�r[VULz>�{��f0�wp�XU-G������qg-�n/vU��'��R��r�N��@	^��s�2[��5^���PC���������h�}l���!��rT!!Q0��Wm�lރ7����S?�A-ѐS�Z��nI���i��
��󌭢�KHw�p��N\"@|e��Ц�Q)jF�p��p�����d#k�-�ֱ�m|��U���:�Rەs�����뀻{�O�� �k�Z��,<�Z�?�Fr1���r\�glDf�ԗ�/�P��z�k.����)�CL���"|@
�9��YM�en3��q�a��_&��z���i���b�������;�M7�턩cx^I�5�y�I�r座�a� Q����=�{���N$�Ϗ@=�؛#���t�i�^F�q#���ۿ�:@ ��I�S� �"SN�Q�����ڃ�E���-�k����6�c�vS���A�N��\(K5�m���C���odg(F��!wjPZw99:}]D�P'3YvS��?ڞ�j���ߟ��4���)L^������r��V�<W�h_��op�wL�ᗵ^�A�T�b���T�s�G7:��ۤ4y�,�����;�q���`�������mw檇U�	��x��%aJ��n�B�XH����n�L��3�*���4P�л��!�ڨ��� 3~E��f�GX�J�!m0��#�C}�5x��b*����wC`2s�D$+� ��A�%������Gޫ'<�"����8j^�F����;?��	��b�v���A^��*�BԖ�K��vӦ��w�BN�)Bp���'*t:f�_��p���� +M�U��x��>3B�d�����tL^M}���%u�K����uszc��d*�+E�� i�?W�pu����;�h�y�h���ird�&_a'�L�>6�� 6S���Q��' ����������|M3

x���,!��p�W��<��VH*g�����ƙ?F��B���p��t�,&���}�.�$��]}D����ԅr�4��(҂js]~5/�
�y�����_7��u���"���횟iB��7ib��,�O���(����������0NYRe���!�^��!�|T�Z���!]�1�F�i�Ҁj�>��y2)���?��E����/�2��\r�z�܊l+A4�����IiJ���� �kx�{��ǹ��#�4����F&֫���1w�3��e��@>���V����`�]kCZ��b�>�n��ỏc�~ݥ�Y��v�A܄6Is�lj����sv�vUڋ����7�ڲ�Z�.����%�����0��R���O�͟�M�J���1��m��ո�J�5�&�>��C�ϗ �rӵN�8g	���`%���B�^ ��k��rHY��.9R��Ęl�e�gu����*�<�&P>���?�Ru�D����z��� �Lq�чk���O�B����3ߗ�q}}8Ȍq���ޅ,�4�����VZ$��΄�)%x-��1_jXi	m���B���t�7����Fo��=�,5NB�J4ɒ�I���_Z�\+e 7&������d�����A?B	i5�I��`�OTl�Cc~��k�Z����WMw�`�&I�D߻�%{��Ω_��w���?���֞iZ>�K���T�@���r�gO}�S��
ꃢ���ͺ'5����g\�[y;��]��� WlS���F��KZ�'�1�J�gf�L"�[�I�

�����p���N?�"5X��aj��A偭��Q �)����)̺�dA��zks¯	�0�ʽ�����0$ȉ��N"Ə�]f���,�ũ��>�w� S��%���n˻���t��-}`|Gj���<� |�L��]W9M��4�����Kg7~�*����yb`ٗ>��0����S�ǉT(y��/gIn'�H�4玟��%T��Z�+s�i�y�jlݭ\���%��fK4�z?������K��v��z-����JZ_Z�,ňю�_��S<{��J�V>�'�������C+�&X���@��h�q�'|w�)y���I�@�c��t���	�3��T.8�BDB~��O�L�#�2�=→k�`�Q+}f	� ���v@	؀�5/��,��*_=a����D^��$���Tj�6��g)N&�M��w,�\���zR Z�KV�;�����xN��ҋH������X�T�M{��sw`��1�lo�%�qZ�,U��o���lDBg!�*������(�{��,�ĄT� ũ���ɱc@O��x�I���?ٵ�
�5a�V7�z�r��w�̷E��.@���ba�p��䴬�N-A��:g���P�v�{��=cֱ��ք-��5�MM�,��$M����&dR�d�MǑ1~�����_Msg�&�]N��V���QwN�$1�H�'>�`nlx	�R�����UT"&�~��#δ�u��Jꚝ_�b]}���}������shz�����FO�*�5Z��̜�3=��_ܲ�f�������/|;t�h�,;�l�T�~=a�.[;��8"���͟�y��#���5#��a��P? NY�Y�K!��'��o�dḮZ���\�Ϊ���/�l���e��R�D���a ���]|��n���u`tH��ʬ�gbJ�tîS�[ѿ�}�Τq?�k�9�y�S�16_��4����ǭ��-~k�LII?���d�*�P��U�P�2��I#f�Ֆ���q�(���M��Xy�՞!�(:i�A�}vS���G'�X�$�0��`���	[ҵ��lgWO�x���d�myu�&͐rX���u-v_	u���������;�V�,�ktߕl[?�S�+�	2���1y*�[@�)��8���c�3qc���aNd>�9�qh}�$zt�?��F����>yu��^�z�@:]��oin���ӬT�~^�$<�#��K(h}2�Gc�������%~�+>�E�$����Ϭ��?H<:�G� �{٤��N#_���m���IX���uF|��R;�����U�[?��ER�Zw����y��[|/V��\5�R0���s)���t�۫� h�� QhB�<7��ZPdK!���[/����~�Yr�ߧ
���@�/oH]�F�l&�K=�)܂|~")?mN=�Id�HV�u=�IK�uQ,�ng����x���mi
��(��[��)EU���_��
�[�!`��D��P����X�*M*�����l�9J�+��ι���k'E���)-���K	�b��	��?KDZp}nIsc�y�V����Q����g8�D-*�;�K�w�aˉ6x��"k2��p/��(9�2���>��3�ΰ�  ��ndvC4��K$����@^R5.��ܭֻ��_qܥm�hE/��'�Y%d��?N��8oA\ɥ;�8{����xb�K���W�%�rҚ������-%��ca^mSD���{���H��n�fⰈ)��"<��[�R���S��P�E��Ì,�­֜�զ�i�n���}�l�H$��L��1�8��GRdWn��a��uR_d!�>�P'��2�vu;�q�:&��?o��[�%��[/��%�_4���ע��%,`zy��X{Ǎ,]�+J&"���U�ʘ`�'���t��ոL��ui7�F�们䟦�xQ�쀯L����JFcU������n�t��� ��f�­ G�|Î�[&s6^н&,�J}����n#8�׷)��,�4(��o�(�����4&���-WD�H�5�&�R$��X�'��e�L�����=Lrs�&��:XS���L�
�N�����u,x^�6��I��SĀa��1'�X�F:M������:�\�>A����&B��Z� ���|@��� 5�!�/^%��\���ɻ�R?ph��w���]��/M�����#��D<b��R�R{����Q���m��A������;i�@�t�>���p4]5.9ϭ9e�������ƨ�D�=�܃������o��B�Wy���.�|LO��:3�p[(8��.���2Q;�����2Y��{�?fYR����y�ܜ�wq�Ɠe�$2`�[nv�vz��e��xx����?>����~P�{���mxE:y#�o���r{wwv�=0��{�f=rwX�5�N<[��LG��B/�!ꬨ���pі��x�/93��Y�'W�ʤ��;�C�I뎄}�a5X����������y*A��r�y�<{�;�1g�T�Ԑ���:�ke�>%���^ {����f�|��/���(�滏��|ڧ���J=Uի�L����} d�Ŷ���_��ag����h���we_���`�<0�`k	>JY���ޔ�DtqR`
��p3��E:4P�7q��P��
X�|���i?��{y����	�hn@V\n֧Δk�l���!���G����D�7͎�B��K���~�W������< f��Y05�t���D2@�e����`ņ���5�|ˈ{�e�v���/f\>����r4�!m����%���ڣ�5����Ԋ�	CH���{n���1�+ePʹ��&�P�����On����~oH_�Ht�	υ����<[�ښ%��j���K|�svk���U�,�^N���`KJ�qi	6�_{��a��c�;A��S�M�s��d!7��66����h����̙�o�e���-����W␏T6�f��;�f�R3�Y`aբ)�0�9#K\� ��glX*�._��:ȱ���)^��}l8E������䏟�,RA���f�&�Q�S汾� �Σ��U��9����	g�-�zc������U^ �;���w���KHݱ�aB�!-��F�|	�Q���C�6K���9S:i�<�_�h�*RzBr�1��{�'�rwn�|�1kA{ i�~^���H�=C��K�wic�eA����-_�����N<;-M����θ����ԁ*�Q��u#k ������ �'�?�H6��o���_�٢:��|��@ذ���ͫ_^0�F�n*��P��G9��T�fz��E�Q�,΍��D�LG1*Qg.�ˉw;F���m�*�"X�V�N���6��-�t�������jU�ϋ�a��5SHj��Q��75{~q�87ް�R�yŐyӡ1� �n���{��0>q�a83l�BS��}��s(�}�2�s��V���A/P�Cfăk�Y����ɨ�ܴ�^���Ъ�[��SF�K>Y�ˤƙ����T�K���/T_��?/IH����������"
�Zwru�(s~�o>#�B�e&�d%�aN���3����4�XoW�[j�w$����C�-�iHG̖�����ƴ�-��/����f��\�֋ wj .~�Z���/сY�e �\���O{�k{谷���ŧ&�r͐u�X&n^s\n������_�"wN>���z>
�|��v��x�UZ}�v��T]}W��9�2h�3s�I����2�Ӝ+�>��*!J�K��?����]�3x��%y��P�9#�K�l�d=s$�H^�8w�e�>Ud�F�3��LCl5�ɨE����X����������tL89r��X�}Z�]ړ�]J����\煈(��Oe6�AX���+���F!��?��п	���t>�jJ8���}�@)��O�NV�S�ғ��.��=[l,���7�36%��G�4d���w"��m!Ų��].�=�ͳ{�I���f�u5xo"�����{ F{������P�f �C/�"H��Q��%�Թ����
\�7��|��h�R3�P�K��o~1�]�)�W3MZ�ҳe�\�K+�wx,O��X�A��gmm�KY�=Sk|�"��2�z�e�ܾ���M-|�SpJо�$P I	���~�����B)���q=��ɑ'n����I�q�æ<����}�G��^�Z��xC�O��a��=��}��^�'"�s�~ay6*֧y^>���܆շ(m����-~]A�+��>�#A̍�5u��_���*�/��w-Dg埠���#=��!�(��m�g,�y������$p�D�^�Hr��=�.tru��Wr��!d&T>�~x��+$��ڟAU�b?�v�6װݐ�E�α7�o��I=����ȩ���@L.�z�xR���y����c�~M6.l�� ЩR�q���[ n,1����H�z�����홣���F!!�c��gR�fmcX�V��r��Ǖo@�w��9��+��S�X�E���m�V�N�5�l�����+��pa�{���=Fa�0i�mV�L߉Gh!%'-Ӆ>J�n�i�q�PڤN�:���NH����I*����x��H��ŹK+�=�����P��4��������ٞ$9���Z�'W�It%�	���6�>�A4�7d�6%�L��5�}J�TW�z���
˥u.m�	ӎ'j�ǀP���o��k�8BAM��F܁�9wٌ`<<��U�H�K ��`�仦�g݈̤�����=u����r����ʒ*�P��kޠ̨��R|�l�i��*ɛ�6��X}d�#��Y��m(8�^�ԷXbI���G�a܅�o"��Qe?:e���@��<p�K8�J��G���	��W�>$�e��8ľW��
j(�v�F*Ո5
�X��^l����%i�&/��6�͉����4[sp_?��+R��2����!<��&��`�BĹ����5���6�ö�q��h�eo%>��wƁD��}��}_����Dg	?Q��_'*�g�Z���Q;t�!�d����Ԏ�h!�1.<ي�7h����1���A̹�68j�Y'H�mhg�\�@��[�z_t��t�9^����6������AF*�j��jr��M��u2�4gOtПA�P)�);�0�ڲ۱�ӏZ'c|�����|lĮ ���Ҭ�'�Շ����&�M$H���d��[���c�����::�*�����?a�6<h��3{��0�b��}~A-���o"r��W�f���0յ~ۀ������k�Lpx���m̌Ld���z~"Y!"�ۦ? ��qT�m�L)�q�{@S��G�����:ey��UF#��dd�Y}j�9�Y~��.N��>�+!�����әaB>���w2������_��-�d�.Ɠ��Ԑ��qH������X����{W�V9ʋr�����aX���^&.�m��h�^zT"��up���b=B��0'�f��32�B��L-�h�}�1B��M���g���ñ.2>/�tN�.�P��Ѫ�kg�$~�u,`}5�.*�u[��Dq�=���\��/�k^��̿�:\Z?�X�
n�u�|���MoN"S!��D�C\��h;sB�=I���8�BІ��1�G0I�:5����.S
J���2���0�2��\��#��q'��xĽO��c�F���C4��/�=��#DW���__XW�Th�-��^D�A[c�F@��@y�_�ĺv}������2Sꊤ*,��`;���Nf#?$�*�+�!=��=��2��%/����h}�X}���0�/i�W��V�57���eB��u�@����A6�E-].��_霰��Q������f��=���H)QGt6����?�����ה<BN�u�ų���˸���(,gP��Y���*[��"�����f���C�	bJS�M�T����k�	Q��YOP��QsEV����|Qsr�=<��eP�y���U�f�롉�c��|_���^����e���Kjs��SH���\L���L���9�����Z-C���Oy�Ѵ�Y� ,+0�mǲxhK��\�3�["y�8��y�;b��7��17o�<r�=O�w��8�O��*}�2co5�s�5ʚ�!�<����ǒ@Az������J��LЁ��������s�� H�&�g)=yVB��h���=(�YI,/��:=?��ƒ�O*#���a���Z��w����+��H;�Ѐ1����4�K���	�&���]��gnbO\�8�~G~������|��]�ύR���8��6�\�!'�~�����נ��>d��V�JL��̬C��
|j����u���`=�t��C ��xW�p�ԭ�v�	��joLj���0���>\���j1o�-P���EF���'��ᄗ�Pa��O�"�&��w�M��kn��ؕ�"��l�p��ciw`�[*+���B��5���5�d7�3�L&�"��4�r�X�%�l�����V2�-.���vc#�[��r�?��ڥ�� ݜ�a��l��2�Y<v��;k���Hl����`�i�;��C�[;���V{�m������Ϸ2�G,��ܪ����4�R���8�P�$���k�!�9�g�)��!����t<���(���i�+%M]"+;�b̗�VY�8Q0�ÞB��㭮�W��mg��ΉSf(�x
&^i���@5�v�:� �A�)2�wje�B��Cճ�2�y���׮\�.��6絛�smѫ�B�c�!r"¥���<,5���X�"���:2:���-�M��(5j{ 3L���c�g$��s@]gpX�z[�>vЁ,uT��VdY~��H��+�$�R����@͒�����I���qʐč⮢���	��HK�x��5\����Ƭ�uaU/<�6/�zݶ�v�wj�&�cխ��X�N��;��3քy|$�0�Վv��+�HBˎkE�'����dte��o�  `����dtA&�+S�X��4,*ܹE<~o*ރ~�H����(@�N��p�x`�Su��g2����Q�8i�Hy�%�G38gƅ�ᐠQEPj��\p�O��/:%���� ��s[�5��Jw�㉔2��
}j�  �Q]NE��f����{�pQ#�;[��A�QѠ/p
�r�9�"BZA��L�LØ�v#⪍7�Q�2�(�y�����ꅌ�]���ތs��g*Y!d7���/�gmTl��� �3���L)6���˝�j+:PzNT�����g�ND/@��a��:0]+��Ajy���(��ӄ��n�p�y��伫pӗ�u��s|]3�I�O2������Q<���o
�]��\�-����rRM�9D���)]� L��h ��ץ@yƐ���q��H�zpi~�󬂛�$m�JЕ�8��W��O�~�*@RȞɗG��_��^{����艬b�����+�~k��>�ni�9���Zd����1#zP�66Op��T3�A��0k;?F��kN�t�'�g���E���Pa��)�͟`&|�Wj����vX�q�(W������tf�F��g4��G2��"7�`:��;�=7�>��=�O���oUMG��j�=kNh���{V��f���	����+%g��5�$Wk��8d��a���$�}B�h�U@2.d-F=�(h[beIcY��؟=����_�qͦ`g�����9��jʅ�1���7f>�5�)c�j�.q��uܩ�&
�Æ�ɣ�V�;���W뉵�����/��u���45q���m|Ґa� �ԇ=7,�&<�\Ϧ2zp,�rK���B��8�3P��K؛&��gxV0z�sq�u�|��e��ҿ#��u��Z�4�Rgs��$�|F��d]���J,�&9��5ns+8�)�0�	�D?f���+�l\�[�(����j!�,��c�
�=|G�C��M�!���#Ɵ��Ƃ��d��jX��R^�//
����s���WȜ��/�O�(�ЃC �\�C���o/� =L� ��ʊn�f"CUS���vn�w��0��O���n��W۸��,OA������?��I�[��lú�͡a~��i�J��~~_u��'��xn8�yd%�p6�_O�5I^��L�r@�-�����}X�7�-�={�o�=���K���l�W���-[ϟY�?������R㋰.�0�n ��� �&���+�i-(�b4�$3������/�c��2�@��=ju\6�mY���]��4ֲ���������t���WE���	�ͦT�Qt��Y�p��� S�����O)���h�4C]V��Cd&�I۽T�|<�z�aH�,�?���~YC^��AmM����MJ8�`�I���A�A!����_1�������fYy�b��J�g�e6�De	���Q�oB�^+R��.�>a� �����r7�`|7�@W㶒MO��&�J�!M~�+��H8I��>��1�����q;�uJ��U_Ʊ�����=�L����C�|�����h$_�>8���-�}��� mY�½õ�fg��޹X6[ll"�/�'|��8	}�^.�y���ȳ����\�~a���|]	�2P��Q���7����hrс}C��̭I���S��ȉ���bb=��P��
�],�Bq�kzPj�Z0�E���W"�]�ɀ�'׎	�_r����DG�_tor6Ըw��^�~�ڃ�!�YxJ)��_�h�u�˭C!�?Fd[��Q�9��K"���:֚9vӤ* <��!r��Uv(��zl������!m�V�J�^&@�x"}�a��$��F�F�k��h�b���}n�j�y��>^;���Q���D�Ė�w�~z��w����8 ������_�lg�1�A�Gx�s���J�`���F��� �Q��Mo宵_�ܿ��ܰ�B�A��n�AZ�.0�g%��l+�|�^!] �(c�Z��7c�,%���88��v�[L���`�7x���5�2^jb�����8�Q
U�N}���;Ut�S�.�5�i0Z��	�(���u�#���D��tg��;�^�6�|K{�jl��y(5͋1nc�Չ�
CH��������N�rNb�*:"���3or�^�e�ԵG֛���������*���9�W��	[x�ז�87�,����
�Ӂ���AK���A�������;�&:%S)����B,�����w�si%Ci�/�wm7�ŶH`$d����Q����S�@`NW$�J���wu�6x�5��a����{����$\�-��Q?���XV�;�M[ÔE��^���)� Q������������m�I�O���sC��RRR���g{3//�p�ef����)wf�D�6Cb$�Ga�`K�,��m+�D�Kv~�X��_E5K�x�u��@�z8N��S�7N����/\����^��9��{l�-���L{.8V/���`�����d�b�����jm)�&�R�o�,�D\yWJ�?ӢđBy�[�̳��tf{="�Kx�OR�6����mL�::A0[��ė��9/ I-��?�Q�{(Tٵ���hB]n�Hnv�,p�V#|���s {9f?���Ŝ�
 �j���-�;~���}k�
SQ���AZ��~��xs�ه��RV�!����c��jD[�K��>%V�A�9������x��B�=p�D"���*��xE�b�RL<3M��t�˗����|>L��ǿI��!Gs�{o+�nrv`��R��/kE���^���A�n_��"�1�11��.ށ��N}�OSw6�e�.�����a	c�,l�u��'蜂<hǠ��A������YT�n�%v�f�$�~˞5����oxik�8 Ҙ�(f|	�U�A�UfS[�}���Bp�� ?�Z�������AGoi3�0w�OJ�I^tkk�6�OxǢa����!��.�BT�׎�pd��5.%g3L��� %��bA*9rn�T�����:fM�tR�ᝌ�`q��!f���ݕ�����\٫ A6�d#�wS������Ng¦�2���L�
\-e���B�b]��cD���Q�No+�HX�;����lG�mDٍdQUCg"�s!�,݈�W�?Z�˸�k��8�ǌ�D�o0?͋f$MgR���='r����{gǸO�B�_�5�mF��(��^<UӖ�gaR�"��?���(}2bM��~��ң*���n�!M�ZSOrzB~��44R�DĐ��P�g��F�nw�.u5 �j��"I7Y(�6���q4f7�-�lg="j	�ퟒk�Z8޹R����	H%� &?�VkWPX�*.$��S���%RW�9 ���6 ak���q��3}��������7�)�������b2!��{�g��jg� U,�.P��Ex��7&���)J��
⨗Pz�,4��~�PY��w(@��D�����>�ˁ���쎤#9Vk0j섭؏��u{�	B{Ni{MTWٿ K� ��oؕ'@��q��6,y!�09 ���|_�uv�߽j�w����%�䬴%7�=�q�)ܗ�3���\Y�͟�r!
���(<'*���r�l}7����D�3���K�l��{��J,DKv���� �0M�e�U;��fꪨ���D�'���8�C�(J:X�Bl c<7GfVS�6����� 6RE5sl�	{O�B�z<�W�i�a���!l̤u8��L����؃�g"��$Y��X"����n���i(Fyz�sv�a�R	�<���6:��/�1�[	`����#��h'���JP����
2'��ĴS����M	��{�'�]��2(�&Q�N=(3<���v*#��4H4Rۿ�ӡMM\h~e:��N���f?��vaT�}�ѶV+r ���M�/�kD^�*A�0�!G<��L`5���dԮ��U��-z&JZ���Ͽ�hg��d
2n`�W\��|oW��� ��ڌ�c#<	����R垄U�����Ⱦh�����;^A�-o-��Hh�D���e�u��4�^�\�}
2���l��MG5���X��xg��[6�_~�"������|����MƗD觖�1��_T.����̄$���-���k^��c$�U�S�]9��rc+�T�>{���>!�Њ���K��t\�fQ�{��H�Z���BB%��0���0�(�~l"f���1@�V}�V�R�Lج�*5�Ar�̦�hTs�Ӛl�S�'Q�|����I�q<D����"�M�-lQ5��1�P�c���Y�WNv�W�,!��ħ1by�\�j�?OI4�ȼ'�����]���zQ�b�.g��5�K
~�d!s/�[�:2���6Ųd���`�O�� O�ynh�-eVI)�w��k�k#9�]����rr��.l�5rI�-��ګq��"�ꂿ�(�۷GV/���Nw`�;mv�y KA�,��~�q�8�w,�ְ�i	**���=>&Tf����D��v�)�=ԜI�ܱE=`����{�*��H��1j�-܈�W	�(�p�(��y)qP�,���p0!�_�9���ldaſ��h<�s������Ͳ�*Ԉ@{1�k:H׮��� w��k�̴���2g�g���:u�~�e�T�5����Q_��X��l'c-���"��Y �Y-6���`�˱A2��D�V���Ö)7��lF��O��.�{����㝼V��z�z���)�5����	��w�x�p��r��d��!J�FB�|.k2��۬E(�R�����n��.ʸ����~=p~h i�r��l,��MT���ֺ��@�eX�x)�~*V_���8Ӧ�_����������*��)T7�.�d�U*�%�B������b��sS6Pu����V �Op�[AJg�D��h&����Չ�'dZ�� ���/Ğn�y��~om��1�lY�U�0 sA������JO��u����g$��2��5S����������j~s�wJ뻍X���M'HDe�W!mnc���A19A��i�|�K�$b��U��,㻍 l>��JK��fM�4�5T�5HP)͒&<{r�}ۢW�,+�b���/�Q�smgu�����+���pDjI���j�����%Y�9�k�|f���0旬25�	���Z�p����uAJ�$�������~J���BӧU��Cۣ"��:�_akB��#έ�*�S̅�21Ytɐ�ĭ�ښ#�8r�t�z�3CmBMw&_�{�b�@"쐔�FX�!s^b��kL�}D�@錽U�A�{�]��� ��w��U�;g���!�bn+��_�z�f�-Cl��B�}!�Q�R��i��픜�¿��F��њL�0�`	zY�[_9�	�$����"�`�"6��A�ݜt����t���Nҭ[;$��Sǩ 2�����:	�W�\�s.����n�����B��o�
�N�ɿk�5�.JkY��ʭ:��~�^L5Ϗ7BU���|��� �7������7�!��{d����]�!�hͶ�^�-_e�x[���L-�g������8B/�L �18VD�KS(Pkʔt��PC�����ָ��$�:z��"�����B�f��>��"尟`}�2e�|��;�L~����5IVn��=]&|T����i���0\�آ���Q��<_�����n�<�pAH�X<�K���&�dxF��ت�\Mh�Na�	x�p���6m�Z��r���S���]߼�
�𥔢����i|X�a"�`q�ެi��rm��ʮb��E��ԯX�# �������+�aI�#���
R1���J(��}��}7BPW�7�?��;Z|%7_�5�2A�m�\��s�x�K&zS��`9��\�r�F��'������D��ZYFpK�Y1�Rz 1�␬R���gIV��|e�q&*�dTӄB��\@�(���+1R0ēG��m?J�F�Y�o��hE>��
�}�'�)Ѡ���ߎ���J#��,�ٮԶ(�g]*�V�9<�A)�*�,L'�����/y�z�&��m�s@E��ڮ���~T����mѨ�t�WR�v�=M<V$�akrR�K���Q3-ӖNJ��G�����EPR��b��O���Aa41�P��h����Ï��Yy�KI��w��$!+_�m��ϯ�Z��%�{�@=me��W#f>����9j��a�
��+L_�ѕ���p�,�9��ք�������bِk��CLauL���{�yŦ�n?TwT�C�҂�xP�?�u�����G��}:2Y#TЇ�2���Ňj��ː�wlX�7��)Ք��[����9-��g���&���m;u��"=U����)N�{�a�`����E��
�C�|���f�h�j���Y`��;��]�RD�P[N���&K������ט�d��C�B1��h�w�[���P@*f|gϴ��S�����+Qt�S�}��Re��<'�JnYpH]��v8�L�iױ��*ԋ��^�V���FW���qɹ�R�Ԋ�ɓ(}a��so��!l;�C�kLf�f���p��x�dB>u��4s�9ٯ����b+�� �nP�:-5��*��bЦeE�٧���f� �� VD"�u8�$����MS�ע�&��D�TӠNQ�f�q4�R+�x*���-��d��ƌw�nzW�����^��?i}I�}v��|&F��ަOI���삻��q�(�^�iE!�F#�
��ǁ*_�3��Y����Qiyo���n����_-�L�iR%;*>�v�zp���W]B�&1�v��q]gh���us�ՙA[HH ����&��]�n܁ewC*uԩf�-�jgn��U�l��G���f�+6vI�=�&��缺���n�6�&ŷ�J���=a��2@e\���6��t�#���Fj��ڼ*T�ۆ�3��ti#�йN��������^nl�fAd�"(���qÊ��2�F�'n`�X���xR�j巁�ߤ�-$�C)^���B�܎�\*��B���_(4���|!�<#*�yJ�⫲�v��<�nsL�pg:H[״�Y��U��?(�UC�X�l��h�N����!iUck���%���+�w	g>\4;R���K�pQoEx�;����_�c����[���S$�p� F�8���h����Q
DB���c^ĩf�ͼ[�HQP~ aU`8\�r]�Ǝޤ`m�@g4 �ׂKt+f͚��X������a�'ػ#G"�4:<�x#�9��\ƀ!#uVvgdd������~��G�w�/��!�e�L�P�� �Ś��`�+���M� �G=�j֝�O#���u� ןKS_�
���;n�4.i��mF��	�62�I2����BХ ���������)�mJ��J�d���8��.?�9-E��Z�rD^��Б9�_�ɔW_�ٟ2�Bx��ƺ��L(ܾ�^�H���=*)&a@�H�0�k�6���y��=u�}HAa!�:�|�h�E��>,�C��~|o�/FI�o���#e}�x|d#�7���]�Z�g%'+\�E�����ɬ���^,}�:em!�|By�EXT� ˚�sK����2��AZ:/���΋����a�7&�9�#��91y��0?���F�i�đ��?Z��^[�I�U	
`VE����uJ-�*�S�W|4L^W:���_j#⼭7�-д���nq�6�<b��r���Wq1�Գ"_H���0+!��F�j��2�l�N����%Ď����d�q`���w[�x��%*d��΅�G�&�D�d~v�T��aq�7餄�臞Fڒ���O)�����y8ڙG����z ����CP��mȴpv%�Tcp�o"k����]��k1ď1��h� ��,�F="Ѷ��}\�I�Zqr��g)G	���^�� S������y�G�`J�!W�12J��t
AJu`��p�����gےx���mb���ϭ��f��ڣ��
��%Wh�@F��`;��^]��|B��FpQh�Y���l���{��eS;������'GF�����A�=�
�B��?䇃�}���g�<L�w@.ʒ��E��p0x,�Ú�]Ҝ�D�ѻ��;��u�w{��k�"4��=jt(JÄ�3?���3�C��4��}�¨���~+bzRZ�Ļ��/`���~���x��E��6��uV��[+��m�@ ��%�9q������%0��Tv�o�Q|J���A#��^=k�C��P��j�2�x���Cz�SHo ����U��(�3�
Hݦ��e��̱�_���ix�'��E�D�g(P"�x�a���W<�����g��͠���:[֎�~��˒���2����S�4;��n;���6:k;F8�3D���Do�Wʝ/�X���Գ4;�T���k��s��6�F��\>~�b�|aw�g���9��T3�39�T�[p��C���pR`����893pN��ߑ����?_�C6���
=���<y)De`H�1ua���<
i��K��BL���0 ?��k��$�^����䋘G��Z�⭰U��������Wި�5�i�x)$��c��;'ِ����*sd	��s�P0ݶ۵���yևþ��n����/�������;���HY�rL}��u��;+1'�6�g��;p\8�.?ߏ�j��\�hL�1j�t~�� E��q3��MDq5���蕐y�6�1�)�������ڐ���u�������fu���z�l���¼���zw�r���g��ɍ���"bk�s�[:Ȏ�-fO��=�v��5�@;Ύ.�r�<��r��~���TMT�͞����Ì�u��q��n�=��w�zÒN?�h��b6�MN���Xok��1$$å��32�/][�-ވqf��;}$��YV����/���+�µ/+A׌��DLΨp4!�Y��tݪ�`tD�m'C�Z��P�T�n�Sz{�zu�#��.K����j$k阷C���@�0�5z?�-�1"�X���f�B��ż��_���-+�$��{C�kz�j�%9oeN3��6F2�"��4�(�1#��zG3�"��d[�[E~��v2I-�Y����L����ф���OkNc�*����K�vw�p[�חO�9�tM�ƲG����s�r�C�\Z:�.9D��c_��Eͩ��vS�
��+���a���{� ֢@,ٌr�!�kT@yA��T0M��%x��1QY�?k����k�>�E��O0�RP���`�!��٦�D�S��Vw�y��jr|^���̕졤f�*��z�-.��fI��o1��J��4\Cb�p]R�}���|Y/H�I����k�n��ZP)���Jꉥb���W5<��	3^�x�q����=�/�`�j�m�<,n|Ps���Q���Z0����a�TX���#Nx��j~&n?<:��C�P�hRk��?�Vc��n���EM?m����?V���`���� =���2v���Aj�q�ml�ʕF�G�}zN� 1�r��~S���{Qx���*��Ÿ�{3\��\h{$>:�!Y�D�%�E?�w��F�,4�4��z"�Pc���1r��;�C��R��$��e�w)�%��8$8"��>����Gs��w��!���>�P�ҋ5��OY[
J	�s�
t��;��WgU=����ޠ��-k�qĺ����-]���\Q�(�&����f�K1�.I�EC%;my�_�͝$���i�X���|�B��v���ƣ�q'����	�n�6��@��C~m߻i}rذ���K�$�%�F:��o���C(�Ӵ�}}��D���Zm�?�XHruV}sؽ =�G��J�jsZHM�]���5'�]�E�y�(�_NX�!f���f_���mj�㼕�:����͙���TĒ�i�����&���C��PT��|,� ���8�w�7�����c�qƬ�ۍ���wl���K�̍�)�Ck��E�O�ӌ`�$ĸ~���zhk�p<�|dUf�2���Y7.�|W��r�#�n [���
:T�&�w#}�fh������H�&�A<�(��T�~2�����s۪&��f+�mU�F2��; ��̌��ژ|� ���H���O<B�͊.��(�6>q�H���S�҃��y����I`�\��IS���rV��O"v���hO*���3~c�>�X!�Xx;���ֆ*6�Y���&�m���o�x	�H��xho���M������+*7>��L^��tFft1K+I	��ҁ�р3���KY(P��fϠ��7�����.�2��Hכ����؂_�� �?,�11vt�U$$�R&~����@�+f]ܶ�F��T�{�u���<?�TJ���tsGa�K#��A�L;rF<K�)�O�P��������R|�1fT���^��{�PL�JY�}����f�����B�9����h9����꾙�j��`k���-X���8��~j���HO���\�K�׉�t�j\ܓ7�����L�2A��aI��F��9<��#�W��q"�u\��R�IɫyE�4Yk����߃��o�Q]Dx���آ�I.����-t���c����j+�(��f��v�M0Zފq�meF�%S��^G�0��O��0]#�mɕ��̷���������m���Z���g�Y���έ0��]��l>j��M�{�8�r!��i_��q�MH��|�h!�0�$���W��u��Vi��kd�E����u�*��T]��%8@I��H��mle^\@�7]ApQϒ�R(�EW_����	�-+J��
�nBm��ɱ��ڧ��?�f��R�( ��eQ2Q	�{�G����-]7z�)�ojD��!�<�N���ȇ��0�7"NC��/�ߚ축�B��^�:��
�2�0�P4�ܹ>���3��`��k%����$�vl&����%K	q�!��a����>���O�j�1�Mpkd��[T�S說KђP9u����_o!��%}��b 7Z�r�U�/���?����0�&X�sf8�iS�a�S�pZ��!�D��t���@q_?�7}oC���;�k%]�"N�v�;���}6<�X��1 ߻)7S�e_!���H v�ks~?@�3����������z�l9AKnI�y]n�y�S��њi�n�8,�i�1n�XK7�y2`�u�%��#�/Q����t6�"{0�h�b���Qd�����33���S[����:\k�ޮOxG�Y��/lQ_�X��W��=�qO߫���ޖ��`0֟C���L`����B�̢p�ex�����2L
u�x��ِˈ4�˰"U_���#��[���as�9��r�(2r���Wu*��4�'�]�y�zȟ��[�)��O�%Y���Yl�v:[�^��_�K���m����_���b�5�T4s}W��W  "H}�y8H�+����qwʈ��n���.����^��$��0ĐtvDns��"��.Ng�l��X�y39��Ԅ�p�S�ᡵ^�u��~Mw�U�8�t4�
�f8O�u4MM\� �w�t��N���Tul�]]�n�'��+�w7s���%y��a���ܕ/�Yeգ�ll��oy�� �#�=�b  rI�*(<S?\_l����}H��w�/V�9�H��C2"2b�)��Ō(��� v�4dy��!+Z'U|}�{��Z�b1��f_�6Z�����S�F|	��p��g���� ����/����\���Л�F�g���+)DYuo��iq&ՃI��Z^���Ǜ�lW!ůU������d��4�"��Z��o��}������Z��������u����.��2��s!��"�Bo�'��6�T�x�P����5�W�`�W��Imv��J��.�\D���L����u��>{����ݘ7u;����j�W��$V��nxWe*��J%_�Ňu��Z��C��/$��)
1×��|"P&�c`-����X�&�2��L #�?+���U���:�E�e��?hn� �	��ˊ�:�1<E�8�8P�n�_�*���cΎtߏ�	a���v�L��&^��y���Z�<_U?��?����G�q��gL"-�ϙ�˓�S4D�\��ڕ��$h÷@��r�h�6]{{��0�%A�i���3��d*�Z��a�=���e%�1�E����X;2�s�b��gOx��9԰z�J+'���=�u"ԑ��K/�xU�,��"����F�2˘s��`SS�	Ј�}Q����ڋ!�*�E��]�H����	�u)GG#g���V^�G��7��
JKE&�'��e�A�./�n�:����n����F2J��Q1�<���A��j��|d�HFB��i��.��]�2��<����繐�>7�X���
�����vd���՞�h�V�e!������߬,ex�k���3��p�Ļ�o���C��ʄ�o������}�/�E,w6+r��G���x��hԽs�եk("��$gIK@�2���'P��8\���r���j%W/=�5��DҶ��]P�eR���T��my�">�*U(�ߣ^��y�g���u9�go���+��i�ٔ;��Q�� h��0����e���sJKj�� p[��A�*Eɴ�[���g9/�(�e���e��^�������M(q�VL�מ��-�SVd\Q�s�.Y=r|��(���ԑZ,�s��[P�S���M���q�/�Q��O��R]�ݾ�:�����j�f)��10�f�9l��~�B�_'�0�J}�ua$��.�bN�H��FJ��i'�$���K�)��l2��Nb5�d�o�ު^E*b��� OsF��7���Z%?o�r�����)�����6���\+�qO-��-��u&�xy�ٝ)Nzf	�)I��5�Vh�'�K�-��^�Ct+^��:t��v"��F"$� ���$h����ڂ��c�]��ٲb:X��=4�B(�=|�G�p�R5��SN��hPN���wĬ2��g�p�Z-w�#TH1�ךr�<��z������m �<Z�Ju�T7~�V��p�a6��{@2�a�G8z���7��c�0�S�n�9//��w��RV�£]��*��j�����F��?�^Ӗ�����u=�-���X�����*��4��ӛW���__�lL�6���W�<3���%�6����F���	� z���#x(��⒙��d�c3p�VH-���Np�����t U< )��M��^�dS���̱u6i������[_��K��v@�[�HN�x��sRߦ �v��vˬ�����bݜ�j�� ��.D�`�9�V��S;"F_q���*���[�X�ㅰ�1L�ǖ��b4��\E21[���Cʦ�L���N��������QW�oɝ������)ZZ�����g۽��.B�}��VO����4���Ax��g=T��o�K���}s �L�&.�fr�1^վ���s��V���:ݴ��\/i=�+_0^rh�h�@ӕ��ʪ�{[��G$k�$���W"qC(��B��L7by�����������FQ�3sȍJ���#-��}���\o������Q[�?��6��E'+�vH��Iz
��k�e��~��*�h�6���f|����Z�Oc����(sc����zD�v�bah�"@�~�ޢ�f'Tn>Q���j���p��ܤ��Osr�~��r\[�jv�N^�"f��C+�J��#���Z-s�"�u'&�L�M�yE�8���P=z��f15aq÷�^�U|�0��u���G����6=�i���r��n`����P���n�*`W�g���ݦ銧���=����ѣ8X��6 K�* �sn�F�+u�ܑ�Q;�T��8~�ږ�<�'��!�݅�a$�7p�x��N�~�0յ>b]���p6:�-_�
z�U)o=����7Z�>E����ՇV͏i��k�
�[<Ǌ��v�Ac�`BCºD|,�>{�4�3'������)u�ǖ0�CZbŞ�%o��ڿ#���ː�a��^�G!A��Ĭ�2%�/m�����A��(�㩢1%����2�F�q.~y�Uu�f�EtBh���������qu9�6&ߑO��*:�}�O�i�J�R�#�0� $%��(c��Ǹ�ӓ�A��73RY]B6=��n��OztOL�Ek��!��ՕO���I��}��H�k��1�N_ǇQ~�L�.q���)!��&M6P�Ǉ*�<����?P�R���{��H����v�	�d:���2 ��\̃P��ʛ���1W�e� �1UGa�����C�g-ƨ'B���#bP܆0�ޯP$^��BL�P�ns��'IZ�<���G�1?��/u�&i*��H(=�G�R��X�lҡ�ݧ��9Lv��\j������x�;�*�fPl,�0�gٚ󔷑�VX�gH���yYaM,���n���S��`�3-��*�p�	/ox,&�܉� и��:�����H��:O��~W��m�����o��g�D�(C�g���n�|�r
�U%�>R�������x�t�|�G��:��(�Z1�%������$ИO�檻��*!�d�U��	b�u��
�[�:`{\ro�&1빷���\;pd��A�E��X��-<���X��R[C�zW�}�7����ѐaJ��V�☢����}�t�5҆����凸� ��h��<r�iӁ=QÕ�s'0R���b*-C`��u�w��]�	�S3���.Z˩9�%��'�����
]Ԝ�I�""�]���Y�t߇:�~�Qu\*\��en�d��]�}�B���b\dr ������y��T� m
��kBd�?5��iF�$a��p���nd�ݹ�D�6��z�ސc�2.a#ko�#�r[�5���l�$"i��>�B�<�h}ʐ�h������^�S���6��r��R��I�*�De���p�'zt�۶9
���?�z^�	��{y��^�-.�&���,rQt�u�v��bXI!x�.���~l��FT;.t3C_u:ڜv�g��I�d8q�^]���9�$Q{o2��N��3���*�c����n�F�QR	1^�Yjs�LY�7O����Z��ēP.f+��f2��[�a����H@cd�1��_վ����}p��k�{.4$�;�׵!I@��Iǒ�<�-Xj���L}�+�s��B=�v��]�4���`�1�������B�����8�<�S��G�M=;��p�t�"��� S��z���pEfQ�hc��r�v��N�]�21|km����΀����ۑ���r���I��D?�63E�., �@���F�Z !�g|���{���~2��z��r!���C�ڨ�@ۜpz/jT��b���TaG���G8��Z�]U�̈Β�G��L�����{h��O�����:���Y�Ċc {E\�3�� gU�x����q�ZR���lp#i��c�t�,�ٮ���i�̅J���\��-���~�Q8@��/az����u�O�(�u�;d�CT��,qv�c�naS�q��T.IV�����-L�4b��ڂ=� q���NO���`�Ǖ�`�߅@�P�`Qm�z��s<����'�;��r;��\$�p
���+{.�����Zu?r�kt�F�KM�^�����7�4� R�μ�{tZ��L{cr��Q^%�l˿�G;nÚ��FɆ�	g?x�!�����?���/����?�s�١�6����$�/	�+[�=��x���{q��/�� AL��;���L��X~(�����R�Y#���_�
4vn�nc֫��c���W�k��.�=�ÒiA}z����Ʋ��JCܽ#h��.�n��F'ֆ�*-�rk&ğ��p�Y��&ǡHU�*H��3��XH8'�.wӂ*���+�=�߿�,ﯓ6oH��.?0��2}�ilC^5��	g��vV��r(�UXd&E���r��g?�?bY�f��S�ё0ֽ=�N�#β������ׯ[(�	��ώ�'S����G�ې%�����X����:
g���T"R��E�g����N��}%�~���8���A%����o�V��{6@�V��|��t��0��fھy+6rds��_ﳯ���OM?^��Qx:��O�lR�����W}�bI�(L����2��Y�i���	"N�l��X�v|=r���L_J��2�>o��c���1q+�� ?�K}٫���Ǒ��{C}�{p��m�.-c�cƸ��qK@@���L���:�aJ����z�[���6"{qd�IO���6�rMJ�6�����P����A���f^O$NB�2�"ʋE�i?�8^j�E�ӿ�Y܆S����s�&�`zn����"}!�uÀ�,r�R�h����Ud`%�x����0x�����f�S<��q�a�$�ō�����aSy���,��ۗ;<X�N@��[��;0�J&{T���μ�޸s5�֊���S�ae Oy)o=Xg;>ӫ��l��9�1�Öv���� ��O��(���<��:;B�P�g~�L<�� (X�D7�׭�劻�����'�5�R��߽w}S�6��t�����^/���(�%��.������6�B��Or�Pi,�՘3h�T,G�ѝ ����������8��L�M��(�[
SD`�/�㗒�����?�Dz^�w��@��õ��Z�=�~�(����<�qLO*՟5����0�C򔮰.�,b����z"��:��.�y���R*��:5�Ȋ���Xx��ȿak�r'u�> koI�c���-���n'.���J���%z&���!����C��3���t~�I6��ۃY�p���0�Ytj��zI�ģ����g��(OoY����{��;UG��\���N ��)����8:1��O���8��Z@��{�Yt)˂F���V�(/���ۙ"���T t���^}�������YY����L���K���Zy�MST���.K���qs�2+>S��.��h`��B�P�?'�J~��GH���l�Y!�
�m�g=D1}�[�)� E%�pѐD�VJ.0� R��Y�_Hجr��8sdR�'��F-��:}�\�ٺu�7��wkw����ʌIu�._�ͱ��Wf��+P��H��yo��+pƤ��$�,���i�Ųm�&���f�.��w��rK�{�.%�2R��˯İ�����
)|�/���\��RS_7�(�BfǞ��f�[G���
Y98�򱼑(Fs�,��^�]u�If�J5M	E�<���4��j7yǄ����w�i|��|��q�ģ���7�B*���*��-�P2��T�XB�ƅDK�m��rn*[]V�](��d$|�"����Q�\���&Tt� ƝB�����"���]��,��ҁ ��T��[ktn!��U�Y��	�S���HD���1���o曊p�9���$G4S:����e	u+�K�>����8��R��鄀��vT߀@�{�چ)C~�T���"b���oC�+���40NA\��Q��tUՏ�5�v]����A�wL�D ��Ղ�xm�L� �b�8"w�yC���`k��a+#K*�:����\�x����5t]�l&W�Hf �+��>�C�LⅣT-��B��Ĕ��f���)h�`�tj����s*����7a����f8{�a-� W�o�?�b��(|�+yLjen��mb��C�pc�1v�mS�5^��*���a2!��[�W�5"�����(F��i����%� �|IVE)�EZ����(*O|�����åH�\'���ҮZ��e9��bSq�^o��
fr��v$�� �0K����R�|�H���ϟAc�r�|���Ɇ�!������u����E�)*�ct�lm����f���@�cN�M$l<�d��L�Sь�T��}�rRp,��9ۚ2����cJ����C*��u��@/�HJ\|(�߄H͚���:iNv�#�xSe|A6�ʘ�QM#�=�\�ZǷ~�{�<o�[$�Z�3�������yS���N1i���_�3e�K���4\��?�f�4�h�;af�w?9N�L��[�˦X��:��G
�y��� / i�c}�=߂�K]G�!��MVu_m*s�PF���;hBo[rj:�V�����\	��DM%j(�C��nb�1�ԓ��M6�;8��p8����Ɓ+>!0�G����%b��tQa�T����f(+cŹ��@�2B�:ڪ�����x+h�,�<�fF<*&8!�.���-g�cg���	�BL��{i퓂�=B���o]vzW"ZiJ'c��CE�q���IH��[�V2��YW��HP�յ���T ��g��j�&g��zs��e*��v S��С�E��f�,e�l�]��c_�-��%��xH���@t �h���!F���X�V�l��cΌ^������Y�q,��O@�g�ǵ��������Q��+_�${��H���?��fb�m}w�(�~Ov��xg��(��Ȉ굽�=��1`�ď���^̆k��jL3E��H�����r:u���A�T�8��k\<Լ_ʉ�ͩ�5A���T�|4#��9/�"i����9�F;�~��4���s�c��ׯ^��c�P�ٚj�N� 4���~����1��,fo�f�p*s䊘j�.�lO�[��i�9WP� 4�����w�Եuw�p�ϔ����;�6�@��x�^��C	s���]@Ļ��N� ;�۵��,5uC���	|��@Dڥ;����̥t� �]���1aHU��P�=e��IΚb5E�J�+@Ϲ�6��K�o
G���-�6�~�l藣�R���w%	�U;����àf|��V<��TS�Z�އmy��C!bk�� Vl�-����Ȳc',�	Ne�a<^V�#7��ΡR���[It�����}���>���P�OW�?fN�H�hw��!4!��fx>X1\X܍f#F8����p�����6�/��Wdf��xT+Kk�x�����7��������6l���so�*�� ;$I%��c*�mh�T�������'�I�.Sq0@!ܬ��A#D�s��8׬����T#�i���L���	Zj��l3�BPL����}�]S'<��¢�A��EZ�,#Z���<q��幙D�����,����w����W��-J1}	TCO�	��eD�b����V�.����.�|�!s'�س����h��Kz���PWV���i�ASn�Ƹ��e@̄�U���T�)�B�������	�!f������Ia������Q�̗#�<k� �YC��b���W��]+Q��Z�m���?�b܄`� ud�Y�o���K�Wq&�
���T���g��`�X�	��ݡ�o�'y,|p6���B�w�m�:'�o5pM.�]vH+Zě���A�ڨ(��9/묔=����T�h���X(]��lV��X�+"bV0F�����h]Df������M3��@�|�`����^,(Mr s�c���ew��S�Mۛ��h�II������0��e芃ٝ�[պbNR�Z�r���@<|�O f�I�#T��IL��� RP��~2fja�.Ii�o��R��e�3j��w?,���h�L��y�M�Ӡ��6\�۱dv�#�ht%�}���#�������G)��k��)���k���,�*m�ٜ�:����]#�/������y��+	�����][����	Br����@�-ޫ-��r,!`Uh��u�7�hxH^j�3��L��x�q4>�(���,�?uЈ�Sf#�@����u[�;F'������ơ4�ia��}����̱ۥ3�t޷�c�O�&��*�?�Ƙ�9�k�1�A��Pkt�F�0Jٔ7���
�ԃ�k����Һ�n���GF��΍O�� �!�uh���%���;���kV�hW���Uգ����ϯ��0�O�6��a�@���*E
%�ջ��V�~��eZ8�Ɉ�7�����p��	���U�=���n����W	b4�8U��M�m^�4�>tcV�DE'�KR�hz���Y��( ����hNJ�$���D��#��M��፩�
�bֺ��e��������	�~�Y�@��2�S�4[_D��GrC��s�Ǵ�P: 4���򓹤�֓�6E1X�r^x`�b-�TAD��O� P=�8�4�Y��#��9���,��z����i����D8*�y�1`T�0��q�w$�<%C
�\1�{���3���Ĕ��<�}x����Q8��8ns@���	����t��l.�u^5ğ���������<�ī
�+�nqL�y�V -�j�׼�Γ��N��/W�ߚG�~{V�uSN�QY��rT���n��}Z��5��J��6}Q��xgv����eKD�
�N����>�n��Fl��g��*���{�5+�=�_��
��B���hE1���UQ�;3�z�uO�v8�]<�]�7E�x=P�����[}|u�g9����l<�GNs��l=U~b��������D6B0�o%uW2�Q�N:(�oI��� �3�r���ǠG��3�Xb�L�w������s�3x��C�TX�&��|�Z_}�����Dڴ�o��r�G���z ��i��<��;�T+��A�b���v<���P	AF)�/��4��&2��7Y!S3����&�ܽ>��$f2F{?�q���y�D��s^^'�ɺUt��|�,:��]��#$�9~�̰>2��r�RJ�ց>Hj�!=~b���
h��Y._����5���V�1����^�M</��E��)tp�+��A�Q���/S�XM�1��t�u�z�)��*{���PooK��v� 3���[R���PNNc�+͋vĥ̐����r!��߭\�U �\gS�����tw$��u7C�;��j<'��������I����W�ư�em�5Z�lΚd(�x���㾑�AU�0v��w!���G���Vت�� �|��^��޹��ד,!�D���Ô��Y���
R=��a��9�bx7����[)��Y�~�2E�!�0+���-����*� �v�B��C^+�ڹ�<H-� +)���W�j�La�S#��kߋ#�&�$�λ|!^�/�},X��f1+����TGx�[/!�ve���%�ek�������.E��qP��@�����u1/İH�3��4�f#*�)%d�+o���$�?�u�����8���e׭���6��L6>9%�J�v:�p��2��85&3�wu�k}��3Sѫ�>��Ӵ�D�֏e���T�	�̚M��'���Y4�F�������C(E�*)��tE�o���~,BO����0��& @:�����9���%���"�$�,�:�
O��[h��'��k�0Z�;��^C�={�h���"y��	֜��ȫ�V�.��vwg���G7�;rƵL�q��ΐ`���
z��$��;.�\�˫��45h��X9�"�M@.6��k���i���sc�e�7xs�qh����4:h�/'��:�,��iӸ�D9C���/�����U�2�П*���߸�l�6�GHRc�^%meM�0�5KGQq��B����uQ11�����C##�h��j������f�\��EH�\HG�m���K%Y�M��g0����]u�^/|l��T^>^�6F#�(�S;\]I$�����Ut5���XzW�5�OŻ�شc�F�w	� mn#�Xa�@M�xش�v���M�T�w��K����Jהm%�t�te�f����<v(y�w�����~�ٙ&��bxH >��� \ƐGR���BOlK��k��
��v���Fc��x���(�Y��d�m�x+�<�xr�9ɖ�-=�{O�i$�ǖ�/t�e��e-����?b)Tz�ξ�f�����V�%�S`�
�F�T�0��>ֽsF��b��X�������@���5��@�Y��:��9p��j�`��*��~���;[�k$�0����I.���ɓ��$���Q�Õr���R�O5��`�?��C:CU�(�Zl\����@�V�m{�	B)�j>����5ˇ.�SR`��ә<%�5،���晙�ц'C�~�4l]��F���X@<��:����;��w���/��^�@lw�K��rj*��/�XnV'���<~���Ά�H,6��J�T;�,[���}׉�ޥ��FӴ��^ޞ����T������n��"�����&�+|��s01}�?>{���ĥY:)��(�A ��U�+��Mڏ�)Y�9YK�]Z�/��h��OwT&��2RM��@(,�}����BH��a �w��U�N���HR`���1���N��E����SI	}R����u�	Bp!ڙ
������\�T\ּ��~p� H���^��:eA� ��B��g�ugv~Da��P�n~�M`���RRx6��iѪ���|��t���\
"��ޏf�wDQm>D�hW� T�L"��xW��R�f�/�4w�B����>Q�뷓E������۹�{���Z�ۄ��i��z�x�����t�'�C��_�Ӈ����gؐ_W4I6�_����S���Ȏ{z?�����PЏ�z�0��`#X_����������������K��o���1�������P�N�n8��8����i�g��^4�Ǫe~?���ۧ����1����?�q�]�%����+B��WgMv�
�n��fk�w�d�-�(NT�_?�����3O��_����B9Y����t?�l-W<\��R���h����(6���ǘ��(n,M� ��g}jG�a6����O��e��%l�y$��s>���y�� 0�_Zz�K��)<�fQ�:��[��⢓7������z>^�~h'j�1�~ OP:$ӈ�#cb�8�WǙ��T�G)-�A‬�Ct�&�C�3��+�Gx�r��ͫ����=��͞�*:aq��xw�V�"/@C2<�
��Ϫ�����?&���8�H����^�D\=�O���-v�]�*y�`N$uO���{�d������� �j|���\i3)T�˛>��f�gT���}�����j�����@�h�eTLu���#��;Y��(4�u5�E�����=��,�B����>��ih�v,�H��j�^R���������\��|L��=:��O��h1�‷�~ä'��ДZ��	������ff��\��*�,d}@k�RcǇ奆7�頉����:�?,�I)
~ǐ�j���p#�<��d�eӦ�Y���P�`@U(`,����W��~$n�#�y��pY2�u:9ғ��������|q�hF�}v�1M�� �.l��>��P�|��8�?�o�>���s�s�{б��y-�".y֦���M'��22�y[!TO���;����0�vR߲~����Jux�ۖᘲPե�[sVւcɒ[i�� 4n-��U;�|JW�\ϻ�g�p��d
�Qf��"IH�)hms�N�c����/���aR���5��iY�-���o9�?�l`�0���T�8��c��Hu��a�K��S�&aS,t��+7ꊴ��,�P�N2���+g#�6�NuS��*9��}�,��	��tӂ���!K�/Qn���8�vBw�nQ�R�k�ӈʬ�k��Ln.�-���� ��9��0$�����f>_��1���:Q�i��k� �h��T��h����]C���i��8iUк8��OcT�=Grk�H�̅S+�L|�97�O����
�9�N����B@ţ��6`u����i�m@0�!�!a�yNТM���c�@�2�7��/���R'��5v35�1��IyC�����rL�L�Y�1Ũc���	L�rB���3A[�����4��yg �H̅�LƁs@���"���|6%�u���@�Q���Ҁ�u�c(�8��$E��yIH�O�m����i��,�ַ���$l��Y�iI�{~��1Gk3҆�}�Y����������iQ~��7�'(�Z��R�w�R����ރ-��;�*-�����knR�|��)�?
�4�V�r�����}Sti��mw����0��*�vI;f����\��
��]H�Y]���GDa����Ō8���%���C� �䔪oO�>�8҄���Or°�z
���e�-��q�Y�;@	ѮV{���%M�U��l�x_���&�!���q�?z4J��C�	3��$W=�S�،���9�)vr��dp9W�����RS�s<n(�K�| {u����~n߀��Z��~7�f��~Q�c^�tz���֛H2(P�	A7�E���-������ą�eUBs�{�S�UQ�C�i����=�����iQv8TVo�����&��͈,����7�X����~�vI�ki�0a���s� o&��ٟ���V-g�L�{{ѝ&��UWZ�+S���gH;��_��{�և�$XC-�a�����iY�l4�b����dᮝ̌4~����C���ϮT]�]���+�$����"2��n�ӛ�5��C}��}�z�.'��N�@aS�3��n�î���c��-,5�!�M�<���R���7P�+�֩����M"F�������ظ�r���}�N�&y��
nuޓ&�����9��7�\	+�R��=�����ob0�瞮��e��rVN|���b�|���ߧb�g-9��l��ᴍ�3T�a�3�G��u&��] �۵Z{`=��ގ��ɘ����NӐ��C��9r�H-!�oU&�Z!�K�:�;H+��D���Z��`�d�IŁ'�N��ʛ�G�����鰉c���*�|�8�i��p�(^0����0��1��.$(���Ӑk�_�m�:j}yR�n�6 �#@������䔲�!)��� i��`\EnK��/��(7�RV�3,s�S�aÕ,��N��tW��j���;��"^#���b����&���K��ݸ�&ۨ� _�����/��JN4�Ӻ 2�}ݧ2�[�}�J����VL˞�Έ�: ^R�r�2�6$.���l�.�WJ�w�[��d��TM�u�H�]6��Jy~0Xn(�c����ƈݧ��� ������4P�_��Ɵw��>����G���6]�)��YũUb��z�8�k#��i��%j`D�!��x~��dMk��{�$0�A�S�ɱl�^*)뤝TF�u}�B�?�����F������Ǌ
[�b�k ����\�dL`:��Ȃ��h�G��z�5�	?�HOqs�)� ]���s��z;��׵/��Ǐձ֢L�&-�ڇd�����mo��^�K2"��3��τVA�>�0+�߇H�+9���y����(b-���n�L�D�����r�䣬��/O�P�c�k١�@ߴSnʔ���7;>q�'D�\�/��8����IoE���5�M)ŷP�3��yY�.Q�)e�e�O�fu�07*���=�6RBז(
-Ҟ2ŋ�=R�[�G��Q�e��DֹH���ƿPG�F+�P�������39@��N�AX�3��VAO�>���n׹�KR��|�١�(�6cX	s{'�F�탵)�J���kq�#U}O�ӱ?GP�*�%�~��2��M�b����^qE������En>�\"ϲkq�>L��wmܿS ���3$l"y�b������j�]S�ܗ�n���i2�>Tx+ؿ�ɍ]]��r�LY�%�����w��ڢL*M2O��?�_�v<��U���CPo��l�s����g�ק H?�j��^�|4XgMq��t�,�]���$�
cs��Z>�c݉��d�������Apb��݇��ɫ�|�� ��p��߿;���ѬKhC�P{Op�-�N�'?8A?�?�xd��`][�Q9���%6K6x�6����m?�|;;���Ki�@yE�;��'���"�7Hj�钕QǱ���6��Z�n�¦] �7���
�Rv'����
:X��X�$���:<R���AX��-�a��9=5���oG3n���i8��$�׫�����މ+���rϩ�����i��N�b�	SO�s�sq���/��X��fݮݳ��<`u@�g
��Q���8^͒a�4G�O�ƿ�������� �U6�`o���ɓq��u���r�a2H,?$z'���΋J�e��*n�!�珅�=	���(jX�>���=�;���˖)�K �X
�Ƕe���o�%W}����f�7�C=i��y���t)��E���L������Dy�p�{���I�u�$�~�I:�/�l���"������~�����%���"�G������ҒR�;��Q5���f 蔠~���X,���h2M�[M�'�w��sX�2�;�"w]ؘ'+H�y�R���� �K�D������w�OD��/���-ٲ�����>经?��z��k�U`������*���}�^��j�������o0Ű����W%[���թY���i����j�:̀�o<����`� I��.�q�D��^'���Ӄ�69��z����~�� 8@�ЖϢ��q��!��?,J�G�G�x��g )tA�z��ҏ���̒�:W���J��љY�O����}�
���y[��\LBz)-���`P=�:�Jg��V�i�����?	��i�},Ȧ�ʽ�G�Lds?U�d�W <,h�O��#��%���h<K�~r��r�#���0"I�a�X8V(J�M���� �DȐ�v�̰�>��w����v�A��h��Eq UT`v����z���+B4D��z.ӿ8����NܬaHJט®��&Kgv'�)v�.|�av�Hc��>b"����o�$K�\�wt?s��ߌ�0n�"�7Ϧ3�Gߎ��ps>�³=}�E���K����5mm����3d���5�"�υ��0խ6�:_gR&�����S-P��	�~�
�]͡]Y�&O!T�Q�EV�L�u��E����\��@�"]u/J^Oy��Y9p^K�5�D�[���ˆ���}>$�3�ݖ&)�۳oK)�6t@x�~�<�$>�z�����	d�J�M\��FD���>�W'�n�����)f�Z����(,�ؽ����2��W�q	����v����m�]Qr)�t����]�F��c�P�o��7�r�TSC���a+2k�d�Y�-��I�_,�ݐR��T?9"e&bS�=myY���J�2{A)9�@�R�@�d	o񂭗�����!��*�֣ ֒!�0��������V	��'IV��0��lN�I�XnïJ��HSG�Gj<kœ�_��
�4w1���`�-�q1+μζ@��}l���_�q�e�i�1G��������H i�B�m)��0[	�}d/U��ƹ�8��-��̘+u���HU,a;j�٩��Zg�!�w�J�.fVn�0c���%�,o�Iwt(¯`��/�'ؘED�k�$�����b�lT�Yo�HZP��	4��7N����
�q	{ۇ��X��Tre�1�r�:�l�=�%�__��-���L���x��):JD6PVa��G9�^V#�L�Å'�Uxe͎��� (��}rr��F"�k�N�@�-m�
�/.j3����Н_kA@x��r�<g�)�{�)&J��j�;�rJt��r�S~YW��Y�����dJ�\(�l{@�oF���'�Ԛ:�����^�QG����f��DS�B	 H]@���Uz ~�!5�K/�և&X���g�Yk���%fݍ\0���s���+��o���Na[9󯹫6���e��&����q�-��_xIքO�i$�dc�KǞ@d� -�{��uL����9RmFhR��ፚu�'�PC�eb;B3���6������K0�ӣ2�FE�Ӎu���G\�E!2P/�߫>�B�P,?���I�*
+�Z�9Oh���vM�/|��h�[5�j`(��f~�C����0�o��-���.1S�X'�_���$�	�XT���nq>u�c�vdy�H�ʚ��-L�b@C�(oԨ=>d�����\�,NyH���-'�f�D�.�Q륲ƫ�類VW�(���ר���Dz��w�J�am������q�.�|[�,:ꘟY~T�X�ys�紏���S��u�q���W?��"�`�V�9��J�jL�'�-^Ɂxxo��pN7ܜ�|#���}���|�)R^�ֲ�wQ�|���dO�$�af���6�Cɚ��y������t¯�^?�.QO�M�:����ñw�z &�&3�~��!*;;��NP�����^�U?N�-\fSP�_0���"��_����Ż� 
�����6\Vp#�p����;��Pb��$�V����`�9xZT7h��M�׉5/�JBi�[�|u[�D<:�'4}���N��_�,"�e]"��ۏ�si���J�
�آX�<�7N%�!SA��4�q�K:�^�#>4����ª�b��M�H��S�O/�Ժf�����p�"�e����	,�_�>/���1�r�S-װ�먮�b� D�QD�b����#}�0�dւ�n7R�(��X0D��s��ݡ�(�<M5�J�H����u��M�2��{a߲���n Ci��~2�tF�*+�"����0{O��t������WLל���q�nokʗ�C5|f�ͪ�ZTV&h�+d 2X5J�/j
�M.Z�E�#�UȚ��Ѯ�T�C)��"�+�~����B	�������� ���┼�(�x٪�_�@�)$j�opq���󷄝kO�ڢ��5��z:�����.7I���JW	�q����v� 0�v�,I�F��ESݛظ\c����3T������B1��6l��D��	��P���G��h�V���:G�)4�--�i2G嫻0�d���W�.��3Gc�Bi��=dɉd�R�θ�*/~n��]Q�W.��\>W���'ش�:#�������u�I��)��AR�{�P��aF�(H|p����~;���Y{�@K0���,��`�E79�<ʇ�~$Z���ʸ�����\Vj���d�!5��hԝ�´��S�s1��s.	���1-���͔-�hhs���^q�����Ȍ�	m��'ð]h-��W�R���o�ؑn�54o� �������s.\���֤�*�-��MD��Hs��Ki�Y�)
n5�kM��bÂ.��u���#�^e����p <eސXo;���u1��B=�D|{#�F����Pd+���ԇ��m�#+�'�����f�gD�5�VL�@�6�e���sc�:�I�دw3jQ�c��ܚ�=-��Îg녰0�4~X��ߊ�Pc�ɸ������T�ޖ�ڍ��3�+�2�h��Qᜥ>TD,�:-�A������� b6�D�+�)�n�S6 $쩝4��lb�
�����:�G���3��pYWJSO�Yѻ�
�"z̋�. �,���������m��;c�^���Q���/�'�o3HNxؙܵM�t�9��N��9�d�%�b��l~D�3W�lЁs��f+�("d��)ua�6Z�h�!\��]�����۹))Q�k���GI*��ڼt�����,j҄)E��@*a�?���E'�O��4=�G��kM�3Q0 �'���;�P%��:̘�H��@�^�������?�UqwhJk�V���p���o�5��q�,.��r�oB�&�w�ED`/��#���xն��g��K$R���D��6T<|~k�$��hv�"jS3;�Y��jJR�qU��a����?t(Wzf�%�(B�U�h�?x�z��y&S���c{�3qi݈^L�׿���
o-��bH�>��`9�yy%J$%W��O�1�=�I��	�����,4��ۘ$~���h�7�C_F7�����N�Rw�5��ji��\�R�6����[���@^�+�}��΢�+���v⹏�OI�^yC�W�qű)PZo�d��r:�׬��X�*��̏�^d�=֦���b`�A!T)�X�*�.�8
��b[�i�%��k'�(��g$-���b�W����C��f(���UU��OA�[�%}�!�1#?�Z�����CL��s�;��� �E���	�Sawuq��ks�Z6-I�ã��#0w��c^<{�W˭��o7�Co&���B)�Ã�F<�<�FJ���{��M럤ځ�S�#w�N�\�@�������1�U|��+w��?����^S���ȴ8 ���xs�R�wsz��{U����l^t
B��C̏����m���Ɓ�A���Bzr��y��b�ru�����u=���?�lȷ�P'�ńߡ[����n$�L���|5p�M����ř�$u�'j�s�ʌ����mK`ӿ��i[#ޒ7}<�q����CbRD�lW�L"@G����f�$p�lYsls���U��l���;���NT�yX9e|�,4�ilj]5V��!ȴ�Z�b\�b�8|�=:�������!̣ǃ�cQ~%��>Y��Lĉ���79��OX o W5{T����!��uO�trҀr�4Q۳P�/�a!'tm������mY�*�)z��wp:X���A���^�MOh����Ǐ�G(�5���{����g�=��'gL4,�,�����e	��r>������g��m鶢\�o��]�z4�،Z px�������xda���/�
�g����*k��+ٍ���o�?�3��o����R<抌�`��w�ف����e��Z+C'�L�;�#4H�#�:oG|��P�~�P
�����U��N4�P
C|�̔�}ਂ���.�o����w���R�v�8��O#8Mu:c?�f7D�-2.����_�#���z�險�? �=��2��9�PV�Yϳ�����W��fE� R#3 ����6~ԯ{���_o�;�>_0k,�r'��pqI{c���}j�^ Ζ�#t�V1��t���ﭠs���<)4?b����u�?^�ѱ�A��hxi���צ�*P,�Fvƕ�s�@��c?c{֒>){mmnD���oH�7���u��uX�q*ܕ1��g�$�a���&��܂j1
��r-���Ƞ���΀+	Yp�3$�8�5w�=Pg���ҵ���fy��C�4��{7m��脫���Ɔ<��
�obb[�~cJE�յ���������m[2������/c��4����������{2|5��ԗ��;��ˠ�K�r�]�\��<��k�բ�D�=OT-L�2�Dh��ł�����㮥�g��ŃΈ��4d8�!e�m,��5(���X�-���go8�DΪE�|�sB�ꇰ#&�#¦��U�`V�r,��F6���қ�>�$������� ��rr����^>� ����1��+١ӂ��[g	�y@[�B�Sf�z�w���@��5����v~r%e�ն}�if�!��y��E��nD� }��Fu�q�VZ�t�\��*4m�D��1�4�d~�qG���U"�5�D�W8o67��c(������
�nW�x}�,�I�.�+%z���S&[��7|�(��K��������a޶���p��=.��fϳ*��D\[ZC8Ci��66�t]�_�7�,�)��z�8:��Vܠ�P�j�	���Ұ�"�5c�+�F��C�wdh��2��ÊNkG��^�)��{��ꇱ�bw��]��.��/�$G;��6ԑ�>C)tN�0�==�B�~�?��8��<2u`R���$ߎ��$NwU)���	��cC��(-%�P�U+�@'<wd�e/^�~���L����O�+/Ր�g���7$-�5�|�Kg��nT����//��GD~T��^��RE�G`��cK�v�G9O��f�*���:�_��"ي��h�zyv$Y ]��㸊�ͫkV�UCa�>�_(���`֡�N����1M�\�����Q�`�|�����Hª��!��n�S����׆�f���ͮ��L)r��L&���l��*���J�"�n�� h�m��^�W<��(<L��]O�fb�Vf3�YZ��_U�&r"�0m�Yk�gL�VF��6�yO	���C�6(��h��a�v�om4�(,<�t�b�0<�p��>8�o:����"��x1����7ׅ��E�sL�Jܒ�іg���\C�%8Vp/ ��>w��Sij�xʼH��M���,�>	�./�`�ɴW��-q2��a�E��u��1���
�UF�6��ҋ�������8�/o�hcbS���6,����m9"��ȿN��ԏ?�(G�2�Ȉ�_��nnXC���9��~�����6bθ�:8��{�9JEb��t�m�*�G~�ptj��`]�"E��1��j�0�K���z@&0n���wM������bX�+Y�.^�$��s��Q#Ĉ�J;y�2�$�d1#d�=|+�Z�烔c�p��'a���g�Ns99&`[(J��LLº=�O���c�����2(��Q܁� e���}�Z3~ ?4r��c1��K�7?]EB���Q��O�w*՜��~�FQ����<�e��a��1RB���ғ�������D�om ���o�ײ҈џ�3�3Y;`�{Ө����TU�Y�s�2� ��X_����*�N1��l9�Exj�`U�&X�j��~ckZA?',>V޶��Mr�gwf��l��A�牌ÍA���ُX�M��TZ`#v�����2/���P�z�h������V=����c�@�6�9�W
�{��۟B�7DX��z:��|�J��ޠ�s�ƪ�:����_�%����G6���,��\l���K�pH2�����f�c��Pم�_��2�+!2�F�	���^�f���Cj�H�N�I������>Z�G;)�?U,�K.�M:0)�.���`�X�lam^� ���)����͙+9`g�,'����8kJG�h�lF��3W��<x�\ V��@eoe<ٕ��`�T�����eo�7�?	����Ԅ��&�".�#}{�̟�ب�q�[��}���-������w�΍�{��E�t}\wy��P1��@x��'_3�^��}�	8��
��LB
4X��5���o�5����J��q��$@��I��!�;�S�S"��y�gn伦>gF@��m�h���~�wɐB�Bx���Tep����K���-%5�X�����fz�Q6ѻI�����Ap�l,c�Nnn6sܢsɓ�Ԥc�ҋ�3��G�9���#�t��(l��c����ه�%�]�W���+_P.ji�]@2�B�^.�S�9�Ō���\�fv2@\�Df��o#�l�qW9u�UM��i��ֽq�W�z���8@*��L����<����z������N
`�����g���^k�RG�sG��Tm��8�C���T ������'��&���Y8� ��D��u�DJ.�`i��ąm�w��_�Ώ����\��j�h]�@�O�1�>,�a�r+�A*^�A1q�>��~>N{�`?5@�o45`<�\�6E3�D�`�Lq~d������Q7P@� �%A^A��=�S�n{ 5Hw��9��뻌�p�Dcv>��f*Ȯ�bu�?�&B���H��(r�r�_�nV�U���4�=iI3���悄d8+�О�{D�uV����.�6׏B� +iPV�u�vY�<����_H	d�����+���H%��A8e�����~�H�f]e�������ɗۊt�:����8?�����  ��];o;�v����o8��w����=Z���N����=a���c������,a�y�������viC�X��M�F�Ag	�9�i�|0��C�x6N�o$��x��7f%^2:�Z��:�6��s!Hax�8,���_w���STyWm�����(5R 3������U�[o���m�݈�i-�_��P�^/G��֋KC��1oehϑZ&cr����sM�R�9�{�>���$��� ��R�v����Ǳ�*�vC�O�7��5�6���y�c�)"-Z�]�˼��$�:'�g˧��8W �M���Rd5�Zϑڛ���|<,z\���_�A'⎱7�>	@�L�#jf��&.��|,���J��?����W[�Vr�+୧Q���K5==�)��E�Ж9��w��9Ts^��X�27�=St��v�'&&�A��*V6G��^s2��fB��CT]��_��Y�Z��_�J����q8<��j�:<!�G�]Ԍ.r��� }d�tN�-E��+��̗N͗e�u�Ji�D/OB���\$p��j0f��]{�F!��D�����Y+�˭a��G���;�ZU�2R�0�U���/�x���.3?��4ѼP/"((��*󱾖Dhw��3��Ee�y%P�&�ֿJ�)�)��qF�_ �$�)�w�E�u�U��t�N���;��՝�ЦZ����wWvm$��&Y�p���ʏ�o��{v NhW���n�E?�� 4�z���+�bl��t6�H�kʴ3��P��H��GZ����jt�����������w}9�E	t�*���NX�=O���nt�	��T���ɹ��Uf�~IU�ɶR�?�|��%��О���9�!�2�5�maI�m\���o��c��*��@�^1��[X�j�-|��<�]��G���?����
����BHt�5��`�
O�p�xR�T�K��+KAy7�M�1��8C���m�a��^!�ӂ��n(�0����"�%x3�u�k�7��{��]��ë�\�<}qϐ^b�vF��bGy�pc8�Z.ب]2M=R�.��j���S�T��7��p��6�s	��w]�+� �xt�!ؑ���z��`��jB���Z�Q5S~��K��P�W�����"�R/�Bʈ�����^+��f2)�jf �����B;��qn�P�D$��f"�pw�K���y�Rm�f�u۫���t[_���
;��D$?�em�ehh	�^(��j�7�`D3��m5I/f���g�̥�L��|0��Mڬ��'�#�&_s�W�'�������$՘��DAD���<o�.�j��LO�Ř�u�����c�ʃ
�]iDtX��,�ʘ~�5�U.6�-�p�g����\�r-{i�$��1��=-%`
���}ӡ7w@���~%qd5@2,�ce�ҨĨv�_t*�nw��TS�Rfd,��J�u�����=����ol8J��^�5�U~�~� 藗�g����y���(B��$���G�b�^��
0��D֨:-��ɴ|��~}��� �;��#���-�)\��[ �s|���$�M��G�x0�Z�#%���'@�-2�ڳ[���;,;0����-�v��E�<|zܺ�|���E�m�z���f��oX}�#�����^�F��#�ه��<�e�V㭔�PG�)w�P�&�j8�cc���
����Cơ]-L��C�	M���o>CcƯ�z��c"am:_0]���N��l&.���U�\�o*&��}`�JL�O�F��X>�W}�a�&r�0��q̗�A)�!i=�܁0	����� �h�'�+N8<"�`ۥ�d������j�6`�D$�^� �w�����J�k��]� iܾh��[�<�t�&��w6��S�8�K|������[�Z[0]���'�E�3C�ᢽ7w�˂L���=���J+�'y�w�}"ҡ;Fp���;��$N��~�+�C�X}�n������!T�9�)d���$��G�H�\ؿxBk��r��m����C�J��R��h�%�:�p�ȥ���G�UM������m�E�k�]�M���ܔ;t�����//YQ�'�T�@]y^DeW��W��*�tQu �9�S|���ٯ�ᙲ &�w�(J��h*�|X8�����c�AN[�|���'zO�h�X�u&�:lR���I��ў*0B<���x�R�o��V����)E��=�E��e�bq˂��ͭНV��4u�Ԟu���� �%�w�Kz4HJh��H�c;ٰΠ����ҵ8�~�π�>��c�,(�ԃ�1Ӹ�T�F3�6�*�FL�^���Dj'�<u�ƽO\���M�F��:�U� @��|��x@h��
�'k^�~��ɏ�����
,E�fU� ���1�zc�P��[�1r~�ƾ���C^d��7ih%���f=Eѯ��]�(�������$T��Ǵ�7�
���E�S��1�q�\�
���h�_��!��ߊ�xY��"5gz�M��##	�N�9�e Ȉ��[#t�u�j1��
��P�,u�^$��WvV��4?�kﬠ����E}��#�*n�(̒I�����߷�V[�Tf!���:���'�A����g �;���%�Q�I����ӕ軘��-f�0$�l~��%)K4��}�f��4+��R�Sr])�r.	Sp�_�oe��l�ݔTݭ�-��S�|`�2H�"!\��a��z��n��v�4��%>�2}���V>TWRYe���>O�~�2"�J&;)����3���n<��ޛ�n�K�?x*-C`%�j��QY�a�b��Q�����-�z(|b+��k�S�L� �KpR��nأߦ��?$�����?�Ύ��O�z�Yp�k�{2t�0y�B���c!�\|�������Á�K����0;��Jm��q��hiKL�������Tl�ڬ�M����/�����U��i�`C�Pя��39�y�mV������2���Ou(�� ��Gt���d���Д)�?aP��d?��Mi���w������L���6˱��.�4w}�o��x|Q*��G��@昿y�n�6��BZU9�l~NZ�ŉW���FТG���Wu1�D|oGzp��͔�����&>�r��^o��yd��j�T�Z��7�������}5A7��z-��yGf�k<j�;w� �c�o�;��X2	��;�`��:p�~#U ���?�u�8�s=4�LV��.S��o���y��o��x�>��)��#�Z\��)4�U��e��|���*�0����~��/�M���)�#8h�+ͯԝx Y�Ͱm�9� �ň��4S
g@7_�G�x�J�.B��q�tHu����>4N��_~����x�� �����DL���IV��QcDC���)�$k���yW���Zo��a�K�����@9D�:�;4"O���Ѷ?ɲ@_r�yn���|r��4���;�c�z�s0�S�3����e�6e�&aF6?�&�P��|�0�<�n�%>n`�uc����lw���M��K$	B\��e ֩p����H��@����`�W-��`P�
O����������*�x�;պ$�E�;}T:]��
+CrSi��M.r:��m.��Q�Ӝi�],���`�Se���R��>r��Α��V�)��nu�5�j��Y������FTN��'�r$B���_R�PUc ��
�Mn9PC^�����Rk��N�`�2�S����j��]Ui�ok+VW��98�k�{G@�C�xv�Gd��$AE��Dpw`\`�C�l[@�{1���e�u��{�bX&Z�Ok+'��TJ�4 f^݀�!��9]=�"��s��84�m6VQ��պ�o}�i�!���{8qK�0��O��bdjժ���tJe�%i��*�C��A��d�1�yk��Z�c�'˙rb=��7;���]�6#����`�һ9lqu*����t1GwY n3t=��)l����-����9z��]U��O߹�����kMFn/�"�I �q{Q*�P���\�$m��� �"�!��V���J<�by�3�liq��d�H�9�y�l��e��Ri�vy��I�톔T�xH� t�Q��m���"r����jk(��'����Z-9�ct��;f�bKR�!5���~U�����wa��#���O�������%>f�z�EC��<�=ko��&N\��df1�@��/�""�6H�Ӟ+A`�D�(��� ���D`P���u8�%�v5Ӳ�+=NV ��꓆oG�5���	�)�E��J�`>[34��h�d�cJ1�R��{�1��@�",5[]���1�)�A�3%2e�*mY�ѠIB��8��mʰ�Ǒx7���[s�Gq�`?)8��5�-��V6VyV��y��b2��f�q/�Ed#+�K Ҽ���v��T��|I��ܑ�Y}JZ�G�^ D�"nҙي���{S������d%KO�ᔶ��e��Ţ��q�H��9��	\�!k>����%
����m��*aLG���t�}�1/z�n@36@���b�|=���B��zbĂ^�����. �����-J�H�8�f�z�ѫS�_+n�-s���I-�!3�#!`ZH��K��y[ѣ�+**��o^��i��z2AX���֬�1�c�-��y�jT�%�+E���#�y�X>��e�N�9�tۮQ�^���)8+�dM1��2$�l.:r��R�K$�SvX���6?UA�a��(��Y��ŝAi��}�ޫn�ͳT5^��ݘn}��
Ѩ`C%[�m�Ԅ���4��s�Ή;w��/�/��`��J���T��H���}���t��Y�+��VhY4h7���E�y�Z	�(��YH�_���L���nX6{d�I3_0���n�N(��jTT��&J�+XLA����-����g ��X�嘄A���Ֆ�x]��X���_~��fE~H8��<���8�oø$e�}���^j��" W0�1*�~�����?K͍�ݔCY�fڍ��Z�I��|O�#0"��"h�	�Mp�ũ��UD�,q-4/;�T�*�����3H�&�p�7ق�+w${���������#Xv4��z{���Y�a{���g9�R�Z���B���VS0���ƪm^�0Mð�������M��5ݵbݱmS�����:Eʄ��͐h��k�aP�q�`�/?Fă�5ӎ"�B_9��)�����
DeS�%�%��
�����ے��8AQ6�9Z�6����*r�*�H����kB�l�:��+�I�O<�s����k�ԅq2���[_8/���X�Kt�&�/��I����h�pDM۳3刜�wüc�!�책��!��D2�y�ķp�٣��;�gV��������e�-��s�N�Q��m3,�����8�J��mT�Nr�|��7ᣲ�N�1p���<�=H[�:�/�QA+���[P�Zo��f[���0�?.PEO�!8��Y��
�ᓅ�q�{J��ps{�#�`\X�����-���&j�����:Y Ӭ6 q���ff��\���	*��Iqֱ�"�T���E����%-����$=듑y�-�	��H�?e�۫ E[�	�i�T��G�����3[�U�W��c�ڐD|���`�ӏ;h�û�k��Sۅe�S��n��~�|�{�{hOgz%�t����6=;���o[���,G��	�5�:��>���o�e
�_#�1/	G&VqgzZ<���Ŋ|���Np��6��h��������H���J�Bӗ�xJ���]Ed�03�*WW��?��
'���f�	ıo�{/�8�	�|6����C5��7{�Sgö���Xy��b�:���1���NC13�xW�j�E*TZ�k�W�F�cp0+mk[��<<6������� ͎�J�<�z� m,2����%����Ρ;.	��̱�*�KQ��=H��`�1|ĭ�p%�'��u�� gz�Rq��k��w��b'�鿑w�G}��kö4AHOG�Jd~���;���/�.��Y�ہ�9|�.�~���0�2����Yc�#�WP�s���/��=�*b�+6�U��ߕ{v�ʸ�M�>4�|3&M1|B��@�+�S�}��-l(���Ri�)h�}��g�����	�U�N72���(�!�s)ì��hp(b���c�L��j��!3S�?��{sP|�ļ�{!��������W���*�@
�U�(��2�ä_�����SML��w{��K{��k�4�s/%df)�.�p����Q�V�θ�g�Z9a�nMӹ�/��_�2�kGL�وm"�U�6��mk��g�7,����F�]�l����q���S˃���e�#?DAn�DȝVg��y��3���i.�ԣG��R������Z������t�a�3�`�`�x|�a��z6+0u�;�(|,J�� ��׍����n��\C�G�K~�BcV�M�X�1P�It����w�rн����[>��E�#]�,������iҧ8S���J:��ԉ��+Y�Ȓnӂ�N_�*@��}mJ<��t��`_��}b���):^���)0��a����w�ˑ�`z��+��\a}�����TA�9��DO�Vhv�z�k����H��#�ښ�(�6��L((�>X(��4�.��+�Ĭf%<�f����^�5X�%��h	�����x�b]��>�s'�ţW����o�+�r4G�ޗ��<m߲��i�ν��T��L��b�_[9Wѡ��qJ}/}�z��<�,�\�[�������=z\���}�	���۟�)������G�%�oQg��A�]Y&�X�oV,i@�����Hu�p��C�4\	�Z��	Q�u�q'z��.ǰu���PY�~߃D�E&��=��BKi�ř����F�W�?� 꾝��I����|��4[��Q4~�4("���`����yF��p����Ҩ|wy����3��P�T24��9d�r����y�B��A`ݿ����sd��}�0p��Hݺ�<!��{w����L�S�L�۔=s[B�f	V1>��~�t�Wp� ]�vD	�J�,�e[�3�g�#�;���2Mv������g��$�?���ݯ:��O����b}lxM�~#��eT�S
K�dDIm(���mD���=s`�5ʐ�㋤Nՙ����k��}��SWAݫ;>��5����2�Z3v8�}��-�~��
�01`��^��G���1�ݽI�#�!E��� �譙OlY�G���[��կ��{��`�I��0kS�K�󕊥ˮz	cD�/}���/��������3`g���L��A-j�0#b�J1u�#���P�GI�^�ϥ�? 4O�L�6ۦ�⣁srdihbЗ�5և��*ڗ*7B�ӳe{��	/�sv{���'��{o�D��=�Z<8C���s�a /!�*�/��|ēIGb�?O��`�C�}!J�H���͐D#RF����Ѱ�9��\�ۈ�!@$�4V�6��$�|�t��̒l��s��n�0�=�"�'��U�L��{�R\��=��99�.���&�����/Pn�������/�K"�7��o�D<�q$RS��i3^I��7�i�D��0�J�����x��"0����5�Q�����z�{(&zB��UQt�k��xע�U�K�"&`#��K�.ơ��m���X�����aL�:>�(N�oߟ�g��}e|y	���9r����n	��x¾�X���x��LH��p�P�­9l�x�=�Ÿ�� �{r����a������䜥�=���镎wLd��㍠����y����Ǹ~�8 G��00����*� ݴ�$��+Ӗ�����ޒQ��9ٷ5�]09�ok���q��� U�ƙ�k�|�f!�Q�����s8s�&R�E>� f�1�"/�(h�n�ޏ��H#�.U��#��͟����{!�*���,-��
�*���3~�,(9^�k�X�ܔ�L^Y1} ���u^o���֑GU:�V,n�?���G��U�A��`֪_1�@�;���B]����
���H��e�c�-Z�!�d`���mrN��b*�ѯh�9쁋y=��g�G�j�\=U"S�פ�ޭ�z���n7q��H�SB�X Bұ�f�n�N�x�6eKT�]����Yb��@�]�H�R��)C)Q��Ek������@?�88s�hU���y5O,jX#�v��u��N��bu[���t!��d�9q
�j��ʕ�`\6�;i�����RY{?�8�7��a�ؑf��TC�VHO�M�]�u	#+�|�F�N��5�\F��e��V���kk�����֣�R��U�J�U�H��\�Rz����J��M~]�u1�Y[/��D\�$v٠�tV��8����)װ	O�yL����4,i��ߪ�1Q�>��$�w����σC ^}#�q��)o�Pp7��+Ӹ�|��L��Rb���L�11Q�~���vqy�W�~�ee`��"Įfb	�����ڹՎE�Ѭ ]��E�����8m}��"���=�F��c�x	š����%�§�1���/o��Q�m��lIb��M�Z�a!��R�+�t%�sE�<�x�2­�a!g��@gw�*q� r��~��q{���#��Џ>�8�W)�߮_�$�O��&.��6�~N�JLj�Q�����n"֥u\�*Q�pc�u+<=�$�� V���bQ�ۭ�_�`���%���sc�Ad��0�˩�\��ʺl���|n|��>�Mnr
/�OjG��*�z�7�cw u\�B^�|ĔHdN��ԯ�����U�Ͽ���xl$�P۸��4P��&�o���������Bccc��z1�6yp�y�D$��?lh����˟���+}�o�)���V�]eܧ���SGj�mV�W[�
�Atl�����L���?_ѕV��9�jb4R+&��t����lZ�x ������-{��p:���DgSU�fA�����(	[R���/$���W[~6�j�9���&�����L
a����h6{�i�Zݗ�ŕD��%|H�c	aLE�RM�e�� 7��_w;�yN���� ���R��)>�2Wmq�	g�u���04���T'���a�B�i�#ۓx3��%DǱ���yC����L����C�� �c��rYn9>h���ow��X� �K�5���uˉ6����;��O�ͯ.���E�����}d�7�P��ӿ���m`�/�ѭ��pL�Uv'^�+=�������骡����>_Y�ݘ�%����{@���z�H��g����Y�������p����}ij��Oa�==��PeI�6����tn|�-J@�;��؍ɏth�R�� =CP���bA���sΏz���"e���� ����B���w�@�.!�|�ۢ7X�>�����z�+�"�zp6,��LBx�G&.�t}�m�[a��P�����g���܈'�9�ǯN�2�{���4D!5b��K��?K���=<�*��Z�J��$Xƻ��&{��&ܘ@:��K�X-l�Q;�������(�0ih��4��|h�i���[GD����'Ø
�g��f��*��$�b�.J]F��L~���)R�\�k�|�ˏf�P�����]���k���(?F��IN�DQ�S.�Ҟ�����j���%F���kCk��������/P�_�s�*r~�U�V7�s�z\.6OH@�@ߟ�ԣ�U�w��E%�pj'��u�q���%!tx���d���L�&���b*k�:\Kַ�c�:�7�ߏt�-۞�=���c�N�ms�~5�oB]�F4z��d��g��:��B6ֺٞ�^���۷�-�(�P������CV7�����+o2���sR�7x䆾u���j�QdoŜG��b D����iU7	����T��Q�%��v��[�V��]b<��7`Ն�z�F�{#�\����&��ر,`���%�$�^�\q�9nP:��k��)�}K��m#J~{�cζC�''5g���S�������$���h��=/�z��hFvBy`L�H�5jV ˷�TRb�;7��k�7�ݮ���mG�'������T[r��ͽJ�z���3GI�a1���N�%��3_�JQF`�>�IE�!�Ew�nZ4I� V�q���\����vnb��(���@3��%���G��7�Җ�]�ԙl�{����Jb5��иKXȢtX3��� ��w^3h8�\ڙV�8v�\��T(�i�-��0�B�I`�3&vVM�{�YC[��mPyN!	\ϏN�U�*Q���͚
�T�Ei�XM�<=^�`E�a���I~M��"H�x+�f�^ƚ[�L���]�
V|�H����%�'��5��50:1l���:��k2򟻝CC��Ȇ���0���:�侫*�q�
�	A�XV��Ƀ����yA�Gɐ*�,T�;��3*�x�9�^�AƯp��;��똖{����J�א�ݒEB�Oy�v|�L�(K6�^W�=->N�k�ݑ_��mj�� �cQ�8 V~*.8��|�T�q/9$��."]-�����m���&�n˓ɏP��e/U�)ӄ)�%�U���(�8z����Z|t&���+ ;P	z���Lj��H��4��X�Ӽh-�iu��e���Һ�����vz<����z�+�9i�c�X��\��S��2���bD�-Q���q<��މ!Tp��%/3GN?��dK�1�!�!|;��w<�h"}��E�$�ή+�JF�^6x�)��@�fy��A�NB���1�,%� ��8��5����WY-�2{q���r�����"H��$[��Gj��`�lwUJ]k?)�-��رa'U�@|�{��"Қ�6�O�䥝C�iN؁O����΢���PzʝLZX�fs�z
��n�`�	�2,���͈_S��5m��+v�m-��E�zZ����;KD����M��� ��rY;e@1q\|�r�)5�{�M�u�_[Jdw�_���3�LQg*J��E]/S_��B�q��ٲ�@e�ş�緈�-0�bX��efC��psP��0�"�'���#��v)�N�ߓ1�s:���&�������-ǲ���`��*��Se�V�WY(��3Onݧ����jt��I��ڮ.9�Z�9�5�9�T���-�x s]>���5
�"�j00����|:�=ײJ��?	�Y�5���Ej��?�{�q�\(���_�S�jy,Q�B;I�8���ite���� �J��]�ʌ@QF�kw���=Q��߈*��'��<>��pvcNt$���ӆ����Yʎ���$�2A�2��ŴV5S�z��lz�C_�o�
ϰ�=�?�F��@��d<�/��~��;�l8�y�\�?2T	w�B+K�4�r|.z:�����/���}B�=m3����L˿���"��Ŋ���:�c��.��ʷ5�u�ka~5,��(��iH�Z.��w��;�D������Z��dpi6a�gX�!�б� �3m���1�ܭ�aɃ�ϣz�Gl�;���@��䷗E��n�V��T�	����A���\!zD����$�Ԅ���[7Q�s����z:N�ؚL<T�/�^)|R
h�Za��7K�+�s�5��Ă�,���y�u�I���r��$��kT���b3�+	@�Nj4�N\}cg|�
x���̕!#���3��rq2h4A
Bm�a =d�ԕeK*m-u�؄
��8%#�k]��N������RO[�͘�����3\Po!s
������z�L �Y
��Y]��n�Ő{�fF��V����c<�c����+�{JT�k�����p&�d�º�Z��^�����_mG�]�Cϐ=��~�qIg3,��eG�y\�2�䴍������M,�7���Հ&@�[�ǲZ��'�Ƿ&����n�ؠ�ӝY�z6I� �>_8���x�����*��~��կ2؋�v�
L���&�V��MҀ+���E�)����L�G�m�Q�����/G}ss�|1Jhʙ�/�\����8z!|��y�c��\lԃD��E!�Hm����1sQ�}9���d�%6��v$�a�f��hNf����Fhs�tf�z ��*��fw���Y�qF+�O��D]W@U��D���?B>4l��,�&f�-F�+�Tz��O��μMz;E�yŽ^�hP����a��s��e����(5Xd�_��%w5r�V�E��R(�����A����1]gs�z���6��Y1��_/+|R�SWNu�|�I1w�Y��#^8,�e'E�ݻ�&���ݗ̝�-�˗�5ML���؅��!^C�h�{����ѭ����r5�����o8������֎�Y��`Ơ�<֧���ܲ�g�T��ݙ6��	C��F��� +\`t��~F�;PK�mL:I�N���SAcN�{�E������mg@B�m�WM2��"����|j]֫�Wp�$�I�Uj�?2�O���k��QiD�l�:`7;�Q92����K�3ZV��i[I�9�!g�=�B똡�7��&!d���y��d[,f�X$� EcI0�*j"�n*:�(�JT*�<�)Z#aI�Ʌ[ϕo���Hۖ&�g��i��ɽw�v���D4u�7�ʔ=��Gh:}A�~�?��\�ˈ;��1���pG:v�OĂ�M��o?�J�M�� ������e�+�H��(ɠy����H/���s#+�4Ƞp��"OI%r	��d�����& ����YT_6ڳ�'<y�Ɋz^�a�'䢮i#L��7�w��qU,I���%��!Vkq�A7j�v�[y���*�^Pk�n�a4�<k��%�&����M�*��Ik7׈�?�.��W}7Gd%�b�9�N�}�&0/7�e��Ueg%��O-�����D�ps�.�)
N}�U	�(J��Q�<�O7p�������$:�+x24�z����ɥW`�L1����{#+$Ɏd�	?Xw�
׻W��!��?��V�x�'�Y8͑E#]"!�u�t#���5p��ju��  �Lf�#a�io2�+�t��^���`&j��H��V�{L�4��%"v��(�խ� �_�>l�w���7��{���J!��n��۫8�{ߙ�1ߌ�~��Q�e�M�����&�׬��?��y2!7�hD'i"�&�BLYݨ��☞~5W���rtu?�U���+�o�	�j �&�k�4z�	�çc?��8E*���-ԋ�"	��`Zeoe���U	��v=KM�x���L�/��U�����Ku������c���o��I�S�S^�޸��>'�8Gj��/I#��?E�Py&���>����(��s�%��x�, ���H�N�z?SmvO� �
������ڙ�88�Z�˦���<V3I���v�)"$�"��	b�º.UΎ'k�����<A�I8I��@��6��}�"��7J�՟r,�I"��U��݄��p2-�/��8ء��%)���*� ���m|�G1Ps�hM*'PE"3��e��ƴtǟ��Z[�,��z	�a�P#�L���(�.�Y�KR�u�S͕1�\����6�3���a&��=^%�~窷R�@
:m����rk�o����?���R��b7�啣u^W�2\���p�B�k��lZQK��X���A-��7dVt�_LC�#�^>�q�ls���,\?�I�W�}��n(�.8qD�Ie��2����`ҟo�R���\f}�5!���j�����3�	���0��XnD[/�k*� 2�}K��y6 aL�=&;D4�1�I��X�	�}4`���jUQ��a
��������o����?#b�r��Y4Ue˗Ad#�/(�.�2HG16*)l.c~#�ڿ� �gS�.XUj�<��=�DR� "�޹���	Z���%Fke�_����wF6��!S5�QP���w,o�8}�_1�<���lܫ���|^ٜ����'Ie jk�w���q�*\��:�4��p�_s�*��`�g/y,�>N��V��ȝhf�/݋g�X�CjO�b8-?2���|e�{�5�r�-��jhjr�����b(��1�v�c7`��\3v�C�G�^�[��������N0΅:�ZO��Q��ɯ!�wqK���eT��9�H�J�ʼ*��	A��x���g�j��oy �X{j�1'2���vi�����p�r�.��+L�˗���lS_1��Qo�������!�	M��59?{p VV���ĩȧѽ�kl��w�Ov�N�xB_�!RP8!�)�k��N�a���9�� P���
}�;��ű�	��]~����ɂv�L7Z��L�q<N��MFe⮧�+��k
��ߓ�;[��G�"�y�l{M!�q)m%��|��:O��J���P�u�o�[*��4�;K�S�G؃BN��oa'o4��%�P�6)�� w��I���Y� (�����������N�t�&��a|@qu���G?��3T��`�+����e��8Z-tm�).UA�;��v����W+>c���:N�-g��v�����>��A�,�+7�����=v�.<�Q����n` �Ï()Z\�Ն`a�@��ț�O�6(j��\&����:$3�(
�}���8���Ms�c%�\��D���~�:�����TjbR�k�ޤFE KS�:^����?��U��+�T�U{�i#��v�2r�@��R;��#h$�Ԫ����`�V�K���~*�o�{HO�՟0�ų��JJ�z��~�����P��-`�4���U�g��Mz�;�ˤ�,��W����ѥ�����ʭ���=S�7�[M߄�"��8-��5�X�X^T��'��;K7�4�~n!{&ut�����!�%��Pv��R}�h&Z�
	�����r��
�<��Lh�N}�NfJn>�+�Վ.C�s�$}&C�@�4�L��p%�1�����FYU%y�����7(T���UM�yB���?lZ7��(�=X��[��������Ҁ[9^���1/�Y�+b͵� �P:N����S!(H�?~9�.���\��C��~)���b[�X��jK�P~c\y`�;h��w�W5~�1 �z"[[��:�փ�I�μ}Z.��E��ɵ�������q�W�_��+�=6Q����8�]�%��
�t���3���VO�&�:��Y盨E��|~�8*(\ܒ��}���?4��.6�~��1i7������=*P=�\���4��p���5����D{�v�\�n���8Џ�<@C^K��ӳ1 ?K&+��T%�b��Xw��3O��p��ד�4[��A���/-q�Z�  �-�D�qO���T_�祕 @�����ዂ�HEy�i�)s���ƧA�ٲ?�"�Dr�Pf�j2=z��d��yf�J�^"�L �Z�%B`2�եq��8��#�$��'h�x����T�E��r0�@\�F7ڳ�O�72�i�׵�Z��l%L&���\͉ PMF%��T�*Χ{*x��[X�5�����0��V�U�,е��o�����4bҖ�~�+o,X��GF�������l%'�[j~�H�=�sz��0���T��w��<V~ۅ�����F��?�~p	`��,|��u&���]n4|Y�R_��2�����(�>0���hD��Nl�̼V�֝�"I�5���E�V�D�o���ӗ�+��4 .=k��!i�$Q�g��xZ�q�V��8^X�����6�[��=՟�s���eU���&�^�'�Q���Q�c��B��J���4b�%��Ϭ�j���4�;��k��t����L���$f�E��D�+U�؝����3��h{y��tւS�D�ࣘG��O�����>V�Rҽ*PU����}��P;��.���Ã"[;E�-S�[��B\��% }�=���Da�[ĩ�k�d��}�ccռ�AcM ��Q1,�E�9q���o���)��%|��)2K��e8���i��FDR�w��^�>!l�/0rK���0��N��i�����ixq�w&b~��C�����x8b�9$G�{����}�jV�s���J�q���D
%��hGN3�Q�O=���+��f+" �`p˅\z.�"�Z�I.�AQ��&K�]O�V-��ß} Sj}!榻���UPm��n�l�,�dX��=N��r����*mO�M�V�LMB(=�U�=!#B�n6e���E���s	7�4�wipGK+��d^5|$~\��ȩ��Sg��>��3��6��!�T-�v|{�����K�}�5$;���,ܰ-ɘ��/��57d���X����
\ꀷ8*39�ü�G~�Qk�O�|�PY��Yu��Z̹��z�5Ҕt��r�θg����� �j%+���p�/�;g���x�_KE$?}�&B�W��m.%��5��+�(f��=õ�$k�tڗm����D�jI�1\,�o��6��C�@��[e K��_�g��۷N��w�x�FJ�����r��˲'�~6�p���#Ԡ�fnc #�_��k	�%���q�gI�<ǂM�S���D�����B�Y-8l� ���+y�ߒ>�:�n����q���,K��S�(�wl�L��}OCp�=�p`]�32k_����c�!��#i��P�����S�	y��fA�����ʄ���hX�8�@�!j�B����a�O�u���mم)�k�&'wT6�Rޱ�w�'B�8�u!ƁM4q��O�B�q](�zſ̨�-�����!��нV�c�J�v�b�4��i���=���d��'����L^�M��}�_�1���r��B�Xϣh��So��7g���	�@�Jp�AI�����?X�ߴ��n�AT�{�Uil���|��zX��`�x�c�̀=jK}�V<St�vhߗ�F�	b=�;n2˝��խ�/[��xb��u�>�S6A��M�hV�$�@�#(�|	�^ ���Q]��3'Y�P��:�=��x���y>��na3S��.���w�.�-���]G�����2T����¦G���mU��~�P����$��T.�A��$�����/�����t��V�ϯU
�~�����f�h�yMU��v:�S1Y�^�g)
�T�u�����mN�b]y��r�b�(R߮Q�4(�=���+�Nȗ�Q�0�v�u�%���ЕU�+r������֗�Gr�Z�u���yr��}�UK
'��d�7q�^K窞��U3������~���eP����84m���/4.Vk#����U_&Zή69��]'ϐS�_���M�7һ����f,�mw���o��	1a���#��%���1������3�6zߐ)��[��_}b�\;%�z�1���7Z�E=�(%��r��f�>�uj��	&�
�*�|��X���M�m�&�5X)�+�K|�:�H�� <�񽋏%��uW��V�۩�~D�M����c�6��*������Q�Ͽ���f:��af����.9�K�0�j~��9(=��*~�����̔�u�,�	����7}r"�D���LҼ��[��f�x	�D��%�i�����~i�������ph2p�Ȍ���a�$�n�8�y�H�M�r���Xu"��Ԑ���4\x%.���[�0�Eʕ�8�����C�����뗽�|���K�}n�� �������]-c8a�w��r�tj���|�P�||���P��Xeb�t�B��Cݞ�٭kyE*��L9|���cL��<K$[Y��f`qD�!n
Nl��F�ϋ�#��~X+�0��a��	JǮ�II�L��-��E�h�w�#�n9��ݏ����Zv�������{�˯��ZL�dQ
7���n����F�:�_�����3&�.��4i`�l?����X���f�'��&K�Ƈ�*@��t�I[n����_�g��˒��G�X&�+{ı�(�� ˠ�n#�ר���\��e���l!��ήe��G:�8�t����'S�� ��RyU/�����;�{�t�J��.�B�P��� �-y�m�� �a^b�~�stuo^�ׁ'\��{�8-I1%�*ܾ� ~�"��,�ǆc�D�!�*H�j6{�ϗL�చU3m	���kB���7���_��4�o�����i��Y�����"������~���ř"WL۸O�\�4�.BB�e�SEH�,��ldr �"���U�G���`-o6�$�%|d�e��j���Cb7��7�6$��ъ�ii�ؾ?μ4}�];�K��
�S��uZ�-���F㠨��A%N�40��36P�8��8�L����8�5�� WK�f[�&^��9�m��u0?1�,hWAo3�L̺'Yؐ��Q7�mN��13 �[���x�I�R�'�Ùm����t��Q��iv�}��L��~��#���h���_��u�'���$����n�`n���D�:�`!���j�>��N�������[AH[;u�����Ĵ�Y���2D��]���b�{M����M��V���%fi��."�h�?;ғz� C��CIm�e���ީ�ܹ�{�v�~�mS�5����o�CW�	�wYM꒾D���F��\�������[�4T��`-n
@׸p�:�i~�	K(�s�U)`D��jY&{x�f�bj�7i�)�ɀqjVr��I|�t�ս���� ;F~�)J�y��/�׊͛p�ꝥ�2m�:����*`��R���9�������
��ע��;67�KH�60BT����Qs�D�"�c�V�� ĲĮ]"�+��C���f;�\M����;�zga2�"�6Ƹ
�3�)~��Ü�^��uA�� �ȅ�����R�Ʃ��7�'y�dq�7��SC�i�~j]��HR�[�P�ioj$.���*8e�=N0>��Y�F�"�����wM��-*�6�\W��W�9_�W�T&(���j�'�{h���˷�K�,o��9*T��Z1?_�D�rT� 8����N�5W�\�Ͽ�@)I���Rjp�[���7v������_	��6�����w�Fr��h�+�b)�|��F��@�3X�	����O�7�)�v��;|���,��D����E6�c|����Gri��^p�M��Ni�j����j���G�Z�Ah~�?b�:�`>�������r��u}���pMZ��>��?�	Уu�n�X�� ��¯ͪ,FY�w,ڐ�:�:���:�x�ت'��MD؟��Y�����aHIf�|WPQ���9m�Qj�֛Hk@"E���OƬ��{ƥR��(X�>O��V1��D��n��k��b��	A���0.�� 1S�3i�y�4��^��+O�*�]0���ä�!�Ws5��!�j݃qET	_������ؿ��Gj�����t=�U#欨�W�u�fA��5l�:zB�/�B���
�~s�7��$�	0-y�Mm�b��v=��s?�ڇ䮑`���9[2?��5Pc��>-��m�:��&_��C�A"�z�O2u�?����^^����dB��A���=	cx"+�H�4��8%������	���������@�	ڈ��q��t�=�YO�i����t$�@�r��as��fZn�!ꩽ���OLI3tyfNok��:���V%�cc�]ӿk!�h�.���d�)��B����Fq���x�} �ÕF�.V���H��K�� ��)ܒt�]�+'��+��`p�\�a��DTڠ]5?a�o�y��H�ӞP0`B�>��
���ʦ��S--Ȁ�E���cXۺL5
	��]8���Wi��v�"�s�{��~/�������$�p3�Ɨ�'����e]γ�U�DE:�fp��}	`�,ό���f���S�����u�q��JI�	�X�X�����­�D��-bEBQ.��P���L�=��e� _��8�z�)t��$f��� k�K(�ـ1�2v(=�ݗ�`8!�^��Έ�C��Ӛmt�W�ؓV����>0��/30b��r�]2%�Z��2�A����1Δ�a��� ��=n�$���t�Bx3`�V"�-xQI��<g �R�Υ0O+G���'�%v�j7��M�J��qt9T`�m��EnK���)p�
���U��r ͂bȅ����ʢě`��v�7U�j���PҀ��1�Nx��Kr'�C�?y����F�v���_'b��'	�Q�d�Pfl�L��O�=�5�$|����ɂ�ښ�������zsʦ�SGE�ޕ8����S�Uy׻W|����^b��G�>5��	N����ݥq�K�G��C�\��6T	KH�<g����l��&8F���!>��OWz]�vB-�y�rY�c����zƶ�ީ�C+j�!���(�N�-pug�����_2,��t/Aj/d�!ݥT�@�f��g�F�3-��~V��9�����v�� ���x���P�t��'���D��Y+��:㶈��HV焖�&�6#�B�A俊Ã�f�h��1B��g2(J��R����~ǥ��H� 0D��s1N.],FZ��o�v%�� ����t9�LN���q���ϕ�NdPc
RJF�L����M6��k�@��4#R3���� 	r�Dp��!��u[^s��uCR��8H
EK���i��[|�{`���P�CO��a�3�2l�gZ'ЩY3�DA\Ըd�,��R�y�W�61����KB�(�I�����(5�{��;Q���@&�OP`o�we�}�3۰��(BsNQ"u����3�KIR��;���.(qGgQw��t�-�;߬�@�b|ˮ)��hu�(Z>`�;G/���TRk��[d9�b b�w��FY��L�SC�M��[c���Ea[#�91��tB�#B���r4D�w�}W�a|n.�ݭ~ ���O�L�7�6g!�3ď�g}�F�f�yJZT�B��=@-��x�H�b1���Q���Mb���Qr�Lj����j?��E.����X��UǗ���-��~x�q��-��|�k�=k�Й�UN�#���b���ނ�{W�xɋr�V�"yq�)������	޽��ۊo�b���f}��,��Ө�|�n-Rp���Vҩ��}��;���b'�����'����,4�>6���~��;2zO`����*����o
��Cr���3�id�J��fl�������Nt�bhU�����Bg�k����]Dh��
qq���R���G�?����@���rH�� <�$�(yNH�c�;�"+�Ǟ0Kp;���'�@Z��\�=~�m#���oh�6Y��r_��H���}s�̿`4]�"�sfK )�]��`��s�\����NԼ�M|qE�$�E7��=�Dk�N�Z/<�����s�N}x`,�[Ѥ�(�� L!zJa�� ����ݔ�r����W�N;Č���*薲i��ӥ��[0|�.�#�� +�!��ʢj��'��m��=5̯L�d��fp��?��p�G����ƕ�Q �����7�����x�Ǻ�cY�]���\�8;��T@����7�>N����x�ӛ�{�]L���.���V���i;����M��n��}t���}�`��Zzߺ��k"����ew=-�Y��n�pl�<!;�!{��1_19�@�� L�Ƃ2.Y@�Ha���L�_
��>�2(B|���6׫�b�iv6GY�� ܀tr,����e��4V�����BS�-�-��C�Y8��@~O?��@t�Nҕ�ΆϨ�'��~����k����Q�����#���R����~���FK�c[�Pj"J~�E-���G96��z�	阀͕ ^9vURU&u��ǮW6�wB\�Z[��{#Q���bH��L���*���i���$즺��/��jS�g�����mi9/��l ��?���]���[{{ LV�>�w� a�B
��ef�r������t�'q6�~�bZ�W.�O�#��8&^Y�ؘ�"�ҟ�^xP~tzkdr��ƻ�]: 9�G����e�i�Ձ �!�`���,����S����*�	P��M�cxG�E7O'</~e� ��q_A�� ��5���+��I�1��wj�����O�I���n�*�,��yڟ��&K؜��G5g�x�+�� ���Z��֮�'�p?���s�9��<�g@R��3;ơe]�T2�%��d���L��w�T���A"b�5�K����vۜ�3�����2����H� �s�U�ўl:q��S�]��<�7GG�Nb6t��f{;��q��.��Hź��N󪾪V���{��r
�#�gת���)���%.4���.�|��U}'�G�v�$"����f�֢9�Φ�R�qէ��X��u�mP�D<������ B��~�;m��A��p��*d�ܾ��b%4�+�]	�3�>�>S�!�#>���$A��3ʐ�N��r�k�5�V5�:�z�d�Y�:��.��ś'{J/UF�J Y:"ӂ��q|��ID.A�������"`�6f��˯�N���`߀�;��O�vaǁr{��Ze) �Vo�W�l�٠��.�nrӴ�z[U��K	���ዎ��+�@�HC���'8�\亅��]�@zG h���"H�VKWi�kg�Ce���pyD)���ް��X�QU�炶Vy��Dݝ9��4ˇ�_����Ӣ�P쐻�NQb
��+�68�tg���]q Q��X;ԲBNc��"�����>�a㚅��Y7(Q��^���v��e��g��E��$�i�9Q�]},��{"�ʩ�*��D�o�d�=��^�-����&�ݝ�S���0̌�7xJ��� z!~�:ǲ�����T&H��	�2Z�ݭ	�?b�)5Mb����w�Za�}��ڬ�>� �yLV]E�� D[T���Y��#'\^��
�ܲ�m�L_ĜNS �o&D��gr3����	b'����S����L��$�Vs��F�s�y�}�U���^�@�I����3WN*ѱ��H�!R�5?lQ����-?׵(�ج�1�܀� �n���$�'	6�2#s�>��������h{���9{�D`\���J���7�F�Q�K��g�H*�ku�����),}8�c���n��L�/>��z9i��O͝��L��'Nc��c�ח�m4H�?����y��:o���~拤f��T����z�0���v�9��BV�s\���0N���O�� �](o}}I|��|U��'���1�լ�upe��<k�f+]�Ɠ���������c�:���� =���v�g�������sS
&�p6���ȳ�ue�����㥋\.�,��
x0�7_Ҹ�|l��\�_n�J���2�@D1�J%3`�� cKC�7Ĉ�᪀��m|�K�'��N����T�i��#!��~��dt���~��p����p]�� ��Y�M����a~lӒ8?r'�߲vZiLVQ�M8"n�Z�4�s�2����:z�yNO@I��@���d��6+�-	��׋�c�j���;أ��	�,v����%t�_5U����Pi�������D:	uH�E����Ä�y�E�����\���6���f66+#��Y^][ �O��*������ �	�1p���Y	y
a��dT�s�_)~����E���m@��W�d9�7kN�Ń*F�ǧ�)n\ՖRv->�t��x��d�MX
�#���o���o��!޿|>�/wI�|�h�ac+�n{ �'v;)�3���A݃�����C�=R9i��k���U=#�>T��1#������H=�_)|x�<G��[<l��u��]] �e��.k���}h)}_d�ɽJz7YzI�߱���Z��ED�I�9p��©?�u�Iz���Z�G��T�l;�k�F'�F���h��Ɲ"�Ҹ�ߵ�!�7�E��h8��}l��9��i�t�7R���)mk���ev]�<�qF|�٢$��7���
�`5���tI�mp�,z�0��]M�$�}�7y��E�tΤ�/�enQ�3�Ѝ�#b>ڽ9�~㈰����>�
��
 ^�'�\�W�֌����'��co�_M��2[�Tz�4����o�&ߌ������6j.����YVm������ ���:�r�;�����l�vca�+m�{��_o���R�tl��ob?T�R��<^�x���]�R�Ldx�y�|"�&'�߱�3�񝝛�H�a�A�9D�m!5	�
�Z��
?uŷ<�,�]mM�e�c�<���q�<r�Uqz(Q�)wb3&Y�{�t+��ʕ@߂@�vi�#h���;��@��l���{66��;�j��8)J�ʾ�bA3᳁��|1sį���"jA�zb��I1���k
j�L!X� ������X��8���sɓ9p�Œ;PC?9Iw��������q�!�5��_��i1T��*B���Q�9��;BY���Ek0mח�C�f�:yk�$���D���.���+)�D���f�0L%lGڕ"��ᒗ��N�:���������nbM- �&�ZH��� ]i�T8]�kt���k�~�c(�#Tl9JV4�bV���.!Y��p�V��f���� |��l58�a��/u�8��M��hvv��I0aRQ��B˯�I��N�T�m�[-=f-V(�6@6�����ڈ�v��FS�-,�\R]���=��|�禝%w�P��jR���9�S8Z-j��nt<�IG���={z���B��R��ݫ�vWG�w����}:t*0�����XHm�>��O�J���
I�R�c����b���ܤ���wf�zV T���C�1��?$ݚMW{6D4�\�6 ����ޕ =h�2ڵ���R)�؅�%�ÂWB��,'��s�30�T9?����X&�l������g\i����	W��`���`Y�'m,��]�6(�����/�����
B�$�/���i{6�m7	���k%(]&�W��-��@�Z��p�џߩPb����̴��#�15]�)Jn�+��.����J��G<���q��d�s�pHh�ʾ��ʠɕؔ������@�Y�Vї�e�����7��N�2o���a���%��<q���u�%[WIG��e���S�Z�:�f��0ï��t�D���\R��ٶ3/���_9#�b=HyF�e��h|.�+ü��"g^&P���Ӵ�1^��{C�_���8�O\L2'JRi��S�fqN��~��Tł:��Md��:��mQ_v�#�*���N�r4��\��O�h�3�D�Y�HӅ�!W��f�9RX=JlQ[����׉����8p��c. `T�h\tl�������/~a�M
�����1o��ꅿsx�pNGա�c�>{�mK����}�c���J-��J两p�oՀ�������[�rVw�����`pD87����ȾiFyRu7C�4H����! ����}�Y�PT�9"��.���S��F�yԆ0��^��ص�a��t���/)d&qa��f|_��éJ�"�>��'0)�T�m^}X�{r��Y<Zg�c�e���߬R��.�����j���G:�l����EI�_-�h�H�j��GK����H���^��6���߀�)���eP��D��!.��3,l���CB����`�%�d;ݺ)b��7'��˥�W�`��\ޝ�>2�fV�K��2���Ӛ5�#��(_�o\ ���pWx��z�����P����2���� �1ߜ_*�ed׌�d|���z����ۙ<r��={��d#T�GQ��I:Iz����|e:�h�_�E�~ড়���粹�;�/�k���*G�V��%�Qr%NI���%�G)�%|�����{D	�~B�x�8%&��\��f,@O��Tz�� M�o�r��yҙ4����Z��ð�1������h�&����@u\�X;j�Sl �?�ݠ�"^�j�ם��Ѧb:9~�4�$�>��:��ݦSvQ�Zq������O�a��"
��[vi��W�o�7�ϷMv��$\��q^�Bu��ʈ�/��(׭Z�*l�&��&�G|� �r���� ��L.�1Y!�d�����}5?�m��;�漹���V�w �,�~�B�L\�������^)�X+w�^��*�ʣM�(�|�a2� ͦ��LL�&ns�T�b�le��\i���G�����s�x!v$�h�RG�(M��:z�\�f�p�*B�p�=,|Cx�[�H�� oT{k�|H
(�G�n�E��I���bV�]Йx`��mb��/����5�_f(v���0�t�:�����9�^�_����:w.�P�������'4���?і�l���	 n�
�3��щ�d<�GѬU�}�mN0'zW�T��.��Z}�����?C�J+�7l�j��pqG��������t)W����n,+~��N�WiUL⃈�p�g���Y�������*���3Gt@6�}�+gy�9��������M��Ī�{C�8U�Y�ĭ�.>pV^y~��9��B�IJ�)������ ,6n�̠�6Q3�4`�����U���î�_>�:�uY��:C��̓|��hG���T&�� �!�Q=9�%e�[8��y�3���/:���\S?q�,٤�˦�`���%���1B�0 �N����
��{8^�egu4�\�{����q=�aˡ��h�S�7d��Ë����k[(V�N �᪍%i���P`v-qJQҸ����%r��E�	FQ��|wK�؊�G�rs�$�N����0DU��PQZ�� b�n 0(:�f����%��ܨ�e����J_�s�����ph��)�O������%�U�����_�n�`[P�jʏH�8��T�@I4��T?����7Fb�k�e!+��Msu�a���຺n��D��';�ʣ�i�GHK4��8��vJ��Ȍ���a�rβ��ww��0N���[n��,�P#�鐑S��λ8�� tX�@؝��q��B���E���B�B��Se�p����R}s&��D�
ךIiJ�R�go�t�X,�>�h��2l��K��o�o5�:�z'7� ��a�~���~@�9��������Ѧ6W=�7�����O����	������X��T���J?���nv�'A�-(��š�i����3�Gw�����t���]�@լE��J�hw,��]��C�_6�f5P�d,��ڊ���XNQ5�9W5��/[!���k�T�䲔0|�I|���W�$e���� ��WIC����� C�����},�R30FGcQ�m3.�M�ޫq���g�}���?�2P�1���D�p -N
=�e]��LȾ>�{ɪnL�7�h;TЛ�3Ջf/�f�.��ĞH��C/k���#p�JL�M�ǋ3� �~k:�ߎˡ�p�]�*&�Yd����H�����6֩3|���" ��o�#����?GӫQ2�#��HY̩I���!Dd(�y��>�f7A�j�C���}�^����\���
�tA�[�t�Zԋ*?��eui�<ie��.a_����a%�|>Mj�9$��b}�_�o��n�iz}�:J��V�������Ŀ�}h���wO���|�;!_GB�'�1�A^ �QJ@<9�<q�w������OSX�u�{��Vא2�R<vXL�\�^�>��V�`_{Hjv(ĺ����b,���i��VS�ؐ��
��/�`�8�����j�����.�.��v�u�TY+��c���*��E+7v�d�R����%ڳ�)�g�����%���Œ)�e�\�u�Ƀ*m�)�Aʶ��Adsg� �Q�Z!u%
	���?���]٥�j�i:�\G�_��m�
��m�=$ʺ7��HE-6�b�`�#����\��(�C�%5�{Lۯ`�	.��
�pW�`S����%����K��x��A���H��C=v�����˖�,���n���3?�&��� �,��$0���k�2'�����t��"�Z����d��*�$�����7�/{=�t�d ����#�K��Z\���XO�N�x�3Q2���$ �٪-���&�UAIy��D~�V��%�w��2����)_�.cy'�Ṉ��e?|?�,��85�<ۗ+i��+t�#�빦H��2RznwE������eX�zr0c����A���J�V��[)$��z��}
rǜ���~�#�M��j������5�FmN�p^�I��0�ވ�偱C��:�c�h�0�:w��#�jVK�H��2���Ʊ]�9�mz:��F�����^	�7�ӆ����c�l����'�3Hij�f�M�ϕa�K���2b�O���\�y!&�i��D�������	!�H�h��S�f�-�7�A��G�����͌)��C7s�v��}��,2�.u[U�r\L��{��BCہ�0��1�&�,�5�J8��ư]IE�'rpӮ������F�����㩄�U�q:����� �'�lB>F�|c^�i`R̲�g/-D��9jOz�25"8����ޤc0��PsN���|d���⡽Ey�Ȭ�t-�Ca^T�'\oV�����A;}m����#����D�υh��d��7���aQeJ_qҥy�^��`b����יq����v���D�T�1�=h82�.@�[�旚z�
�t�廙H9�?�E�(�N�*;��b��P���^���T	zو�Eh�6�8u�9�㧨u���*����O�\�:�k���������L��f+�Z먞l�m%>�5����kW�g�F�ǳ���[iJ�kЃ�'
��0V��4��$f�W�X�(���n|E(�~�F5����R��̖���N!��O~����&�?$�����C��P��h(
x\i
�V:�~���6�z����'���,t�?�Z��v:{s��ⴿ�[�Wq�,�L��z���������pZ��R�*����J�L���i#y����o	u]�vⶽ��BM}�I�a�D#��{������m�4c����?A�ϸ�"#W�6z�+�}�!��q�P�@�|�j\�r����8�������=h��>��3�"io6�G��Ӷ�_�L��̕.�;����/��zt���4�%�"�Z�5�'2؄1���n��%vUIl�2�����,,�"V��RQ�>5 �.�b��-��Nz01�l��bKfz�6Z�Y�YQ�we�6(q-I��U�P��W��3��G��.��@m���7P>�X�������;���Ñ�\D�
O�*vU����k��>�AUc�h���7]�BM0�?"4LA`�l&
�?��qs[$f����ws�W1��>eM�f�������p�C�G�����:= �*�*�r�~�M�7vʀ���W���Z~��%����.��: ���_uqh)���[��K�0G�ǉ���	�"���U���ˏ�*���7+"�c�҈����>�\�Q�! i�<
�s�^y�a�]^�z
�죔�D��#����y�?��'�D����<��dcJZ$Su�D��J�@M�$���v��I:ߐh��e"����(�E�V�B����t���?�>(T�����k*��b��O�nL�
D�!����G�UY����p���W��"	T�#�����s�~��Py�:5nOfX���~����G�����&��.�jqUH��E@��"���n��L��Oy5�g�&{W�T���*�(Ɉ�Wl[���`E/pԅy�m��p�;��!/�AD�����8�Hf
�]D�Ϛ�Km�qv(^+2D[	��r1,7��g��M���Ù%���\%��T٩'2�"/���ΤQ���=�m�����x���1�>�;�AF6� =�kz��z;�~L��c�i��<�8�X�	wn��l.wo}D���<�J��i�~e��@�|�k e��cv��0d��p���q���}g	ڔ3@80[�ϝ~zD2���rKp���Tl�@�� ܭ_<��ظc��^��bJ�����859F�ί���ZI��r�*���j���b&�&�/��`���h����d�><.|)v���2��E/�|�\�5:����A�m�2�bfy	*�~��8iL8�@�k �Eh��tI��@��I����������������
����g{�~�Jأab�c�&]�K�d6�`e�l ���骟���m��N�����	��L����[�Yk"��o.h*��:~�g@k�Z���e�N�Nn�Ti�Ĕۥx�:��LihU����Ϻ�`\�p�������O�z�͔����S��@���!�)��Y�v%A�;�i�1��\)c���	(@:rS���:wH��6���2QKHX��s�g�A����gp	�z����H[�9<BI�) ������كS����wm�a�	�)hb:DrM��WU�t�n�z���g�J�I�K"�m�S�с��h���Xi\���M*K�=������� r�f��U��*�.��WI&�Ͽ+F��`r�l��#�
i�Ǩ:����-�e�u�}�a��Ho��C��F�rQ�{����s6K�aꘇ<A��{V궛�[����C��T�9v���,8X�v���pwu1SϑHR���9٦��,���蜴����Bg��fl�$���.�F����1(�e���ۤ��V�Z0 ����j����>�~�b8�z�Ra'O�
�1�r}�\x�SU7h�Ƒ���F^"_��,�f���T�$O���N�d�Wo(�	�rӂ-��MQ3�R ���H�I��Ҵ�6R��M�a]՝CP����c�ۿ,˻��ֻ6ۘ[_�~D,�
�,4�
�$����ï���y��O��1*,-�{(Nra`�K�κ�lZ2ɿ�!�fd��6᧭ٶ)�S��A���6
S��MT洭�i!��uڴ��-�޿0LMJv�~G�_:�$���b3#�\�ؖ�T��ތ<��k~�̎X*�O-�,\���F�'�o=�5��2�=,�%Ӿ �F���`
�W\�^�U������.�l7�ZFk �Sc/�~��&����#�1�y�^�	!��SGy�C8f��*����*m�=<�ܥ����H�X/C��r�[��8�x���m\����^�ޖ��&7�y�����ϗm�W�|ݚ{���ܣ� <���m�6�&Y��Z��l�#Rf}�B�����*��{ 4��Vm9��!M+/q����(�f����{�\�/_���M���*����$fp�xn�EC�ܺ~���/T�B�|��fm�&Xh� ���ݒS�f�C~Xu)��E<r��.��>DQA:wf���k���i�j?a)���B���tAs��-���px���Ej�EZl��7
�\ii�Ҍ����g�;�-��.�\��Y:�T��H�.��[M'�6�����i�QzYKH��Rܦ���@:���f�I��®Ms@�E�����+Y�5�mT����Z���:�π�s_�[���'F�.��pv��Ըa| $��k�ÿ݉Mof-��&�^>S�S�d��w���g�9;^��l��@>?�0������x�2��I�#�k��}�.�P�|����w�ieS���[��gN��"uR���&���xxI�R>�Y�p]�7�P����~[|��n-�ُ9�4跽�>�Ģ� �
^��"�_��	<Ȁ�t�~ެ^���6�*\
����*l�縵�m�Y������h)I>�|eL]y��kQ������q�c&,O|%P�AG�6��xq9�����P�KJ�ݽ(ˀOPzH��n@��uܰh���Ї1B���?z�Z?r��%a�RCw�Ԙ�$e
)|}���$7������1����w�H���2�#k��=j�5��նxm����x��H^@c{��@Gǟ-#mX�q�=("���~�fgGȔa=�\4�6�Qk���^it���L��_������윣{�����^s��C���rlz�1Y6�VF��e��1/D�a0�g�1~	��dz2x`�)�EA��ʄ��C��Y�l5���
	�����[��B�*H����5�=̤�G�k)�:=��~>�̈�8ʟ����X�6?]��0c�`�\�_m��B�ˇ+)�'���xf���'������{�� ���W�r|.X��z~�W�#(���<�P�mnlm�8�#~�<���N'#g_��M�٣�z\ԋ�y�\]/$��>�g��hMS|WC$�F���?�0������|�G&�-���*.�\����ޛ-�n��4�I0v����lǇT�����-f�."���mH��A�<���,���a=h���\�� k���.��X�Hۯ��h���]�A^��>4zũ���l��U��̹�i����Z��б�C_�_2O���~��'Tm�BE��(�7���z��o�u4e;,�\Ə��P�[G�?hi�h_���Yޑx��!;ZNJ����P�k��绡��?y�ŋ}<d��`��NU�>(�������z��ݾ�@=�-���Ժy{���<l=�FF�k"�ETXW�\�tqSr��D����N:h}��AO��Z�%{u�Y���������\��@L���Bo(��&����Z/h&�ҼC��e��8��U��2���7�IP�Fiο�ER��ΰ�b���LR#��LU~)��
�8U-	�BWV
�D�w�r��[�������-���9�f#D:��m�UKZX�R#-8�뺻]:Y���ɩ~�91�	��)D������(�yM��Tt��}V�������}����kJ}�/�y��KRԋ�s9��քD6Y *���c߷D��G�w�~������Z�m<��b�O���q;�GB̚��+�L1XJ��_ʺ@�m<�w]P��4:pMkiw�m�#�96�}@�w��#�;�����U�PN˟�AÝ������mB,�8>[U��Ӧl+b�S%O���4���Jt���z`��ggu|z�E��!R�ZMlpx�r�i�q*N��[�A���?hg>q-?=Z���~i�D�ܜ�$Q�U�#����R�����k��������S���h�;� 1����d����M[kdD���t�h�������h�m��G $��\]�;*�_�-���B���ҏyx>C��S���М�$5vA�����g����M[��ڜx������F�(ǉ��k��%	�i��b����5�*��R%�Ы8�X��4(��`ҽ�'K�O_Y��i�?m��|}T֩P��`s#]b�bj�l�~�ε ��D��p�Nh��S7H��k�' ;J좐o������N�D���<�/hVJ�n�5��W���$��&,_ �8G�F��t�@$ʽP����&���֙��ڌ�o�&%��^���l<P%q�Y�P
W�]����ê�oH)�U=?�7|.���R�]��⹢��Ck`�T-�DW��$�#m�NC�%�����2�r.߉�B�􇸚	�$:Yh5��H/I�-�ψ'!ܖ �2�8�&ns�����0�D~�Hp'��E�.�27�
7��>H���2gw�_�)��3���33�w���mL$�e�Y��rT�c\�����i?�9S�Ƿav<zR��N��x߃	W��Ht����[�P$�U�4�a\�4'���K��5�U��&��z�H�c�t���+�A*`����./��6R�4�7� �6ܛZ���m���r�6�܈�rR�ԕ��!�+�:�kJˢ�_7��53B�[K��YFK�Ê��(;DO~�M��AK��s����>}�$Ym� �#H����!M�����]u���\О�*g�0�s-�	��vy\a��4O�z��֬����=�>}��|%�a��ե�'�d)^��B�g����!ejA�/X2�4盠_��sI`�tL�����s�l,�!h����ly�x��ck��a� &���?���7:}+���ĽSQc�>�t���PFE��+ʭo��@�1�:h��	#��� 1��L��C��ן<��%����	����\u<��M�t'Ի�v<(�~�RK`����Z<î�T���(<�/��!?=�����ƃ�7*	!�?�uN���d�w����3�����.�����;��M�{1f�xV3l���E���*�N�S��x���CB_�Un���P�k�������<\�ۜ)�?�(r��#1���o:.v�RM+��2�u'n����DMtH���B��u����D�0��<��+��(T�m�sj��6������6��P؋���.�;��I����9����k}r\� uݎ��ɼ��$���v��χi(���VjU�@&�0t��k�C�d9��6�
.F�YdD���@(��~�9��1����s�y)q�c��À�����R2�a��3�{�A��Ͳ���<�ZM�x�]I8�(vg�b����N
]x��o�
2�vx�ݔc�*�$�p�u%3�)���ΦL���T�~K�N��Z>v��vv���L�p"��?���rȡ>(G� -���ʔ�Ԧ��.ۛe�~;DidaP�;�#�����&��~���]Kѩ�ϣYr4�Z�����Y�m ���5��"Χ8�K!Oא��4]�)'C*Xo���:��2;e��|u�:�O6���^�v�e�υ��un���6P��կ�5�i6I6��������j�1����4��1\��:�S��8��T|�u�������1U)K�iǅ�upo;�O�E�� ��`�P���O(6(�W��Н�C�9a~F3�k!��&�:jA�s �V,�:cщ�m+3���� V-C����]g�R�h����,`P�����b�[�',��/d�.�e>S�7�7>��E�Bh�.30�D,�JÝLg�s��pU����VQ�P.�,�g��Y��cr�%��Ps{Q$��G��0����x��à���2�GQ`q�ֹ7N��\� ���o�]4Ok Ho���:s��5J%�b߅o:�e����53�+ѩ����yK!^dI�EW�xTHz�Z(wxMp@[��}��@ !I�ӡ*�2-��[p49_d�L���-";y7D7���]$�������'�	��z��4�$�;�zc��=�\�
g&F̖^���z����G�3Y����qU�_	�]"���<B�^_ҵ����+�eo����)�0�iA=yA?���~�w�WS!�Q��ek�!����W�n�|A������i�֚��?/�%'�nj}MUt����9�d;�y׻�C��(���@/y�.7�qM#ʭ�B#Pe��Beأ�)�};M�&�6�F(Z~��Ʋ��A�ҜQ.O���ӯ�*9k�Y���?��l��X��&N�d��H���Tb�1�N^M`��>A
t����%�
�P���a�'��r�G��W�w�8�ii�~v�K0na�MT����1��zlY�H��r����Gz����n�w]ȋ5��i@x�}��b���5��Ѐ9J�,e���w���CRj-v!��曅��WN���^qTZWw ��J�ِ���� pv2�,2Ϳ��h�X�.$�(q�� 2�����!=��N=Ky)�'���c@u>�f��ɉEWWq�Ȳ�$z�Y����L���u�L��vD�,Q�!��0�#���/!�G��ݱ����r�h~���Y|\m	��~l��>B���[k�ܭ�3�����6��1g�A����N�Ď�O}�a�g�'�4�U��?�
k�����wc@&�m91��%�r���/����wd�h��� ZF"�w����ғ�N�RK�.�l�����<��n�T�h['C0��ΥL���%N�V m�/�Y�~�r�q�131��s���Оө Q!$L�Ę KH��l�1�\*=�m\ $�Z�ta�K��S�G~
�I��J�ۏ�
ݷ��s{���L��4[�+QH΁����O�i�x�Z�k��7�%�W9�g�KŦQ��*n�ɟ�?qp'�'r쇫�fО���ip�nj���&ڙ�����RxJ�yV���5i���~��u{�-���ÚBO��mX���O��UyDu{4q���1�-��AK(:��E����"q���4Dt5":����� aeޤ|��]�"��~@��˥QVbul������̿46�*�h��B9�$��5���>�#GʯP���Οn����ˑ�Rp�GM�sX�ٔǖGz��D����v'�ˤ���T.�b������[!��zvT5Tr��`SZJ+`�:���%�u~ ��k�>2Z�\�%ى�Q)�x��g
�c
�l�O4��|�tI�m�\�P����Say�����f��yM�ObFl�.'\\F�/\α�;��d�&@�EN�k(c�"P�y"JPLOC8�$zS�̅]���� **"�.C[���ln�\���D"��q]>u��^`o�������w'�#ىp;�H��/ރ<�&d�yG 2V�T���G�(�C3�&d( c��?��-=U	��0��"�c���Ķ��4��n>�6���� "��/y}wQU(��S�w�[�L�+��)s�c�m�Vg�%�e�aUk��Q�
b��g�Fy\�t�s�n<�fo /O ��}_v�,��q�˷��E��^ʠ3���{v�Q��7~,��F��N,B\��!����@��T�U�A{�O{FL@����oU�L�w�0�i�Ҝ_&��F��r�nEy��>�b�E�����~�9[���(ǬX}.���؂Z.,SP0�/+|�����{Й]��j[��^Υ�ܖ�f��%ρ5v��V�i�H�|v��ڐ�}�����A�wė��S���Z�vcvZh�������K'#�����O�)8�ٕ� Kl���C��2&�O�I���U�c�K18����zDһdF>h^��#!�����!��vq�ս�C~3�u�OiCr�2�66���ѥa����|yo'F�pp*B�J��#��׸U���p�]::;��}���+� @W�.z���L?�,��"�AV�FJ�\l����4��c桎����i h���'s�C^8w��$��M���a��u1���-r�:R��ED�[���	��eeE�&(�
�<����m��DC�1!�ܩ�Q�bW^��]���+��m�|�uŞ�ܢ
��V�I�P��s"��Ʃx�R���nK��WJ���8�*^�ȩ��<�=��X��>ɺ`����!DW�fvdIY�~oB�/X�V	��:�RX��Q�������6��͞�>Y�=�%%��]^6�%�4��#�.�a��7��⻤&h��ϺX$G�ĝ�֒�2Z�dm���G�����-i��R�U����k#4!������k-�,06H�����mO��5���{����쁴��응�ԪSJ�<��>k�O"�i֣bҢN�3@ ��b[���K��"l��%�|[T�������y�f�k�cڼ.7W[ּ�)��� �L�=���2���c=\s�e-v��sf%�=Vgb6+"���+���M���8��7y���T��7�v�4��x�ȥ����+3��'�ڊ�"��]���,C������ܟz�`����ϲ������V���F��90�l�Zh��M���@��ݶ<zVH�M�D��Q=G���ǹn����7�z�G5xwyP�/��C95�q��<�
޼ �f�����TP��x=�#���t22Օx�I'���b�C��:;���q�EOHb�.y���)]�K:��SVz��k��o�}����o��s��[�a~��<BL�1�3�X5@�\�!z�[�hRK�B���:�6�h�}fK������X�	0C���]eg�e��\��kz��ABA�ј�0?f������/���@'�x0�(\����Zh�%*x�%�9c3�!_٬�>�dk{���z����AѮ�͏��()d�~�9r
���g��m�ؙc��B�_�"�p�f)v[�ASh:��B����Y}� ��䉃�����1#Zf��yn�C���r�R �z����t�×u�n1�I��_�BT�ɟ��;��<� �݊�UG�u&Z��jrtT�����D`
�]���ҕ�N8��ng���4i`:0e	��U����x�d��+Pj?1�s�����J�>��C��k<���7�Æ
��'*��4T��o���(%����+�H�&����0��	�<[F��眔f�#�A���k�l�LPɚ�pl
�o��&'�^�������k����,�����Soh~�o�t����)�n���|�yu�9s�%M��[ܣ�L���j��sIӲ\��$u6��|�y|�����)\����"���$�c�B���9��%�2C��.-�d�.w,4�%�B��*~���`nڛCk�B�瀿W��n5-�C�����j�)��9���d�AR�DFFĩC�R,}���_k��S/�1��3uz.��]cj_����O#y���O�Ax��������ڶ�HG+����pnGB�<y�=�<RK�O�f��t�m�ˢ�A)�� ��N��_O1��8��q�E���q�ԣ895�7hfxb{"�0?���z��*5z�o�t�����OX�C��"F �U�N��f����Jh�n����>�E���I�s\�B�������:��X�d�!*�D��_-&�~N?���¨�f�ҽ:�L�/�!z�w��O d�K�&a@ 4w
��?Thu��ӫ�6���)�/<4KH���]�I�?�ί6��C(���,���ha:�x�����������z|�
��k��p6�g[���'�j�+S��F���w] Ν�$����8_»R%�_�֞�^)+�oP��n�� 1�*��gpL�}9@�%�l�°�*M9�b���v�2h#$��  �<0rO���yg%�D���	:�#:����g�hEĵ�x��;�������.��o3F�[��W������y�LѾM�;�g�+\3�������oO�S�1<���x���*D-h�J~e\�N�������w��������N.1������B S�XQe<Q��SMpM�@���;G
���>���kK�Eg�yR�8�	���_3�gw��'T�f~i_l�u (�ſ":ڌe�=�~��@��LĘ�f5ib.�W0��A�8�{����Kk� Z��[S�E*�vm�T����C�������%�
�Ӷ�p���l&<����1R���B��}�$z��J�j���e=:�$!���;�@G�o<O��c�/���CW�>7�mn��s@z�=l
 K��|x%�T����:�S�����ﴎ�T`ґ�~�om��2����Z�?O��n��b;߄��o�'iD��o����	�Ojc1d�T��El���^��:����a^�io=4[���އ��A<�_Gkt�g3�Ҩ��P��O�k�#�D����LS�ȗj������ڿ�6�n��,��̛b�X4$�Y8�tޟ���j	�q�xP��B�W���8��@�Օ
u����%q�޿�1 ��Y��,��7��f��������<V�0�j�Ƿ�~?Kn[�l�¨QUH7`�. g'Lk�]�\͎�[��ۊ��зU�5ggr�6M�.r0���đ$0��y�o��ܭ�c��!Dq���\#^�'Ũ���ІL6&'��������[*��_kV��\o��W�(��gr�$�G(];�q'`ހ�s�jٗ�%�G�S݉lυG�_��������YH��jV X�����lf���ʖa
��ժ-۷�J@n���%Q�fk,ߙ�����e+<����\� ����✘��U$)j[��#20/V��`D�r���KFI�<�M�t�IRUѳ6g[ML49֍;yoǤ�|@څn��M[�@�G�(��i�H~���Kq(���]2}+�������t>�wʌ�9`��
�	��r�R.�	n	��b .V�t�kpėd��O��\O>}>�m���f�j�K���%�O��F��������;���W���X���P8��)a�٨���M�6�3�d�S���ST����w��Jr���'3���b�~m�ďŐ{�N`m����w�S��t�1���hӰ��=u#�.Ib��������`a�:G��k���bo��X�!������!���=�i j�i�A	C��࿜Y7�ƭ1�4D����'bW��2������Q��A6>LX��m��� M�Ջea���+{x��n��46�}-ۓ��G���k�q؏Yqԗj@ ?�1;�M��2=������%�N��w��_�3>��*����>6;�<���	�4k��n�p|�ta�S��u%�ѵp��j�U�����>YZ���9�E�����]&"�SL��g��[��p�x�d��,�ٴyd���cɚ�z��}q8kY��̣B�p�F7�����?F��� ���9�W`�8���"�奔<�~$�SH�86�G�k��sDG����ɥ�����*��vd�XW��
.y��>������̚�l)q���1g6
:<S�I%��	��0׳�u�x�uoJ����K��뵰I�R�H~0��>���w�*�� ��գ-�d%��Xe�,�_bd��'J���vجÖ��8�G����-x��u�N�9���&NVU���ά�"�Uߠ�ص����:�|�����o%��f��O�j�	��2��D=C��[�r��2?f*R`0U�l��נs�!��S ��dQ������i�5,��u��j���0�cL�3�z�n���6,M�V�d���?�rC��C�\�^�I7�D�Dqv"a�w�W�7���ڃ(D�W8�L��Oo������O�noS��;��^�B#�h���p��>=|JΎڋUk͋*���3
�rwB	N��V�H���)B���l�䧎9����8/�c��[hz�49�=BScA�iR,LM�J�!V��3l����alBW�P�T�WMl��yTRGҊ��R|���Sv���M
�s�� 9%q}�7�x��-��eہ�2�dl�I:D��W=�H�\�~�!��u�f�B' jճl�pS^2��lnY�����1��i���a�NHo�&��<��q�n���$�+$^RI��:h�*ǭ�@�I���@���^:z��Ë.*�'�_	�6�"�!X��e� ��i�r��-��ëE�'㿯<n7�7Vf�*@LN�Fd�L���r׫<d��p.��ї~����X1A�,T�}/|����R�tX	7k���N'��2��O�^���*~Ww1��҃����"�n�������̎����^�5�;&�y)na�(�_�� ��@yK}�Hbn�^�RkŚ�Q�&��v��Ú/u�ʽl��S@���M��1̔��j��_���l�u/�o3G8X�w5�W��Wj[�m?ɞ���C��@��	���<��h��FMD�U��}��Kxۙ��KJ��#�&6�?�Ps��f����Y@�w �7Z�*#�wQ?���4�~ߺ�H�����z��_Y��8r�`5����n*!��һ���-�%�]��:K (�������u9:1
��t���;{�CL�^�d�f���j=�2wc|���3vx.�RF/��ڗ�Z�r�_"�=_$��Y��o�I���)C�^G�7Ƨzܛ��"F��ֲ��R�5'y�r���W��hA�X^��q�=�:��5��KC�(��k}�.�{^�>ɬGf����3ر�s�uU吿��ũ0:�5��C�g5���{�����\o1�,�|9���BB%�.�F�����ﳙ�׳\"b��L�Ǌ2��\����Y�sR�]'�����R��AE�V����~z��7}�Ae���sb_������g�2��Fۻ�EB��-�W�<�C��j���W�8R �xW4�����.6�0�L�ͥ�lJ�g/� T��y�3R�>��xH�?~�)�<��q��b��tw��t�Y?o���S��5��ʂ�r`Џ�1]g��Emt�}R����?K�Bi|5מ�L��*r�V���<5ݧ���In� ��-�X��}���e���D�|�{�.h�ɔ�5F�|�[su���UD�$d����l�Z��+�3i6/���j�뿴 I��˴�>���m��k-��_�|�O.�e����0怷Qˋ���~��͈�(�o!a�*@�CwSQg��U���=
�P�.2����6���m<�Υ�o6�X7'��A�vह�6�ZP��0�.�e�𗅻��:7���D�,{�$Ī^�j�"iF�^l� �����6�ήK���A�x����O'~UQȐ<B�I��6��(y�;bT��'\?X�ωC�� ��Z�d9��+����Q�f�R�hǍ)o X�xXC�w7!4N-�4#nz��p\�X�PP����vgQN������r�J�"w�]o�nq��o�+%�3_��!'�`�i���	Fg��5�^�$��p��+'1/�w�H���(ƙ��Ne��>d��朄��B�< ������xpo����Bl���5>�TG�?s�O/�:A��gyC�v	����$j��yo����i	f/��p��ټ�[�ϛ�D<�i=�f�99{C9��R����C��?�|�61�Ȯ��N'��Ғ9����k���w�3s���ҁ1ϲ,��u���ּ����9Eb�{�~�*����[�(�dñ㑍ci�M�CXS�n�����?����`��QE���?��V��p�鋻C9?��C2YO��|��ʻ��ܶl�̺����$�2zѳ��u���$.�0�K�޲3.)^b��Y�0I${*����1j|���=����=�xcx��e �̝�IÀ`B��-�;X+%��}� ����u{p�X����I����n^�)ZG[�M��$@?��uW4�������C��:��m�N���1`�t��w��]�~�_4�%<�Ә�'#'��N} 튞&�U��O+����ڻ2��  ۏ�&�N����Q�	���Y:w���d���F��bF^�X#�t,7����T��fV�Dj�����D��o���'R)e��2�O�W�xj�[gQ�%(�i�@O���+�x�b�z˄�;��K�¼�_�_"<��%N7���̘x� Nu&���Jd�N\��Pܩ�&ܻ`���;�<�^)��}�IT�}�a�n�El�����i�4V���r~u���˲����9�Ԣ~�{X�
�?}T���Tԇ�#����n��5x��$��R��ҫϯo�1�SZ���\��P	5���B���]Ѿ��h�%���d������
�r��|?���Ao������+��������7��<�
e��&-��]�s�X��m7�nN0��:��I^)�2��ՂTޔ)C[Y�9J�b�=Zd�Ȟ[�n�w�	ln� CB!$��AYV+��]x���,^�g��\j T�mka?�a�����\�~�m#ELN�RQLT}��CE"ת$��`��(b�n^G��$��&eJ
�P�3���k�c�fP�7bCӆ�I=�p������ ,7����C��4_e����jO�/r�9�\f��"�󄡏�^%�� �b]n��.�2�朗��D�����<K)�A��<�K�l�������
+��dL��˪伹����v:�B.��qA:q�v� �@ߓc�n�m���S/��[�$xe5� /q%�f�=OH������	�kw��]�.��07����-�%J;��`E@ھc��+V�3z�uD�zѐĵC�����T�e��� Љ��%�xr��L�;�	� l�U):`E#T2�=����о�	-�u�]�v
:"f�uakBa�AtŠ]0q�&�l��V;�������Q�n�K!�A�c� y����Eό!B�T��\��u�]����&��b��g���("K�&�?�O���(]De��TX��\��4e��SP)�2���T	��Xlj}�e�F�F 1���	Fqp5x�[ˮ�k���2�#���6� l[4�j.v������| ����J�{8��R7�q���7�t���
'�k�2�T�Cj	�%�_����@������q�+��n6�z�Z�e��Qy1N4l���_8�.�aJLp�o�agY3��s$@Vf@*��hF���XLx/s�"��
�T$�B8N0?�!!�h��%ѹd��|0延qCm��
p���5�_)�a@[7���ߙ� �7g�i���O����N���˵|�^���2~�h�d'K��:@f,�a�����m)d��H'���)-I��	�'�q]����8ե��fi�v��
,(��<?��$9���H���zs	j�i�c�L���,�����Ϥ_�9Za}R�)عdtM�'�-�W���Ѷ�[=c�%Q9d�SA������g�����`ہ|.��v��8���$Y���M��y[eT�a �=b�
=L���ۣ`ޚ��������z������������0��2���$�&�'�B*1�� �ǣ�'w�#���	��;}i��t����ݝ���d�QA9�	��I	8�H?oR��DLͣ|���Xh�g?�k���v>_=H���{��n��(�����절����܄�~�a(�GOZ�����eu��VG�Tӝ���.�^n'�Qiś/�'؄9eF�t�c�lC��>I��r g��$?� �%�{�L�\�av[�t���3sT^N,i���j,Ɦ_��`v��o$lC�{ѧ�-�pWGù~B�i�{��̕�K�Pp��iG�8>�6z����oa��zk��ϋ�;�o�(�I�%�z�ap��۠~-�B��m!:x��
;��8�Z��[�l�Yt�F6.Ep�!mr�N�|�~�C�ݯ&#۲��Ɏ��]aMQ4����áХ[r�3�h�a�����A��BnR�θŤ#"$R���j�f0u!o�@	Bk��9�h����.����x�Yi3���v=����<qw	�T���bP�8t�+YJ���bY	x�����_iq~�+��Q�4��P}�����ct�� a»���`WSζꔮ�e�K]�ͽ�������`0���(�1lq�(T�������5߃�H�N�l	t	��]F�0������RVE��9A/\@/�B1Wni\+hD��U�0��eήލ�	/G@SPS�it~D�r�B� �}���Xs�aǑϟk1�a�i����&�O��5w<�-�b|��>3)�5`�s)�jV�kf�F.�8{�X�b�
t+���w���aD`��������NiR�'W���q��T����T�S�c;v���F�w�����<Ww��"��,xz,��*,��qb!������Zc��
K�)�!\������#�E I��t�R�b���|A+~��.�e�)��	�H�e���>�l��Ҁ�Gh�0��#�A�3�m��H�?�M#�`���#�z��'�rS>��2��%�,�m����?�Xp͖@�e���@*�a�K?�
�@�^�X+��M��<��(��G���M�>��q��'<T�mm\���j\ى�o�4�jY�:�w\ ������HBAX&�Ȍ/>��58E��)�C����.zi�yN̂)��([�zg1<ż�,3�[K�9)	�T{�� �U(�O���;��������[�d���]���.��-�νq�z����芬q�m�?_��˞#Y�NDO�]��?r%��h&.ڑ�kN���+�4ˇ�<�+u����a!�F��ZH)$����x���B?���Q�/2�2�*7R�wƒ+@��^�h�3G�ֈ_�M~����]c��o����9�@L9��z\u����r����#I��q��Iy�5���xZ��W�n:�ּ��p�yVnU��f�nu�Aw�i�
u�K��b�"�9� ��~oa���1��>�d�\��y� y�3́r� �S�����&�����yD����b�K�$H��w�s�ē�?-���XD����8_=��d_��B���J�:fI��].NL�J�j��֌�1�­8�y�˗���t�t�/䝁�a^��H�Rt�2L���f����[~���\�q�ꠈ%���\���s����ٓfk��|����Hj0�H�������{���n�������Q�+J�� 	� �����N
�yH�ǐ��)�T�J{���g!��?�H9M�Y�� �0����׬(��3�[�ޒYrZ�k���SV}��&1Zo�>"#�i������ТҠ�;[�I�����*|�Y��s��/���;ǗGy5F���u��:��D����Yc�̀,���"�Tz����s����l��l�z.�%�u�9��p7��J) $���=� �'�V����.���O$h�N΂���J�����.L��dDO� U/b���VnǮUD>��*"P����73�'���e#lڠ�U�~W��'��߯)B?��<�!|-�>�5h�ٯ�e�3��@���=�@�L�Xz�of�Ń�g���]������(�4��3��n)��֛+G�#�FEW@����[gOM�cs�����A8�-�*:< FJ@��_p~�s�/�G�;�
�������)��-�ULuS&���K��>Wg�!��R@	.s�S�x��N]Y��{��H�R�W�]�(븒���[r��o�|o�� ��J�H��ωH*��	���f�P������%��L�L�YO춼E�o��nA����4Yl&� ��/W��׸{�UI�$�EA��٪v�O[V����p(���1e��I�^n���#��E���+Xw �r��p�qȺڕ��7�4M��|Q�T�V��Mb��)�%yʝ
&FO�+������N��F�)g��j�_s(��u�3�<y��'���g�T=;9����-�Ý����Ę䁃4@C����+zf[��[��^f6	��2P�Y{���z+�(��
���N��޲g��k��~0����=YC�]XCsu����o�5����BA�����g`+~�՜H�6���.@�̈́I_��cy�[m��!�G���M��Y�*
WC�(GѮAQg~<^[�E\ro��?y8��`�.��Q�"��u��%�����hBK���!ر*<��!ǐΩlmFc�T�4�-�3�G�%g�X�Հ�f���yϩ�H�g�_�=|C�6#Qנ&
</����	����S�ZyP��85��t@ j}x`!4K0�i*z�}�q�G���4�������5d Z�~�����KJjĥ��6)���E^粮 �����y��6�����*e:���C$�U�R� q�8��Z��f�Tq�<!����m<M��!.��U�&@�x�3� z#��&�.볯��sfƵIM�Y*�G��
錥ϕ����S@��A�ċ��V���N�h�H3��@ Oq�_��Z�E].x��h�b<R���_��C·}*���`��1G���]={���zف��3�UMF��A�5L���z�9���c#.R��ا�A�Œ��w`��o�7���)� 7���2B�SlЂ����=+����[�ȞEJ�A��MT��$B\�J�-b4Æ�?�9�9M��˩ؓ�����g�_9�sK.
���Р�@�{�OS�]�pG�U-F�h@�qo� Px�K�Y�}D;�\�2�F�`�ٓDN� �=-�XA�x�%#Mzj�Ʀ8�p�k[b$�+y�:Ì�3z�3z�[�9D]y�Vm�p�4�ҋ�8�=Lً$_��&B��§ ^����z*#.�������?,1��ؚK��%,ַ�Z���.��e;�ܒ�U=����g�θ =�a�]"[/�Fb"�[�pZi���P�*�rt'��`g�I�}��$�L|��R*1Ҩ�9TFkvǴLy��X,�y�'�����EKh6�M˥'8`�ɢrt^!Ow�"���4;�u�kj�����~|�=�� M��ߚ`���3�aW�h-sXi{6��F������
�^�*�!?6&��q�J�������Jz�;]�$q���zt��.S2kk0��h��YD���G�|�ނ�T����gZ�����h�����"��O�	�����q��y��B�g\�Yq�����cY�q�LX\MI�US�c��8@:���%'L�����e ��F������νf8�����C��3���&%�m@u}�T���arۊ��s�ӹ��j!� �BIģ�}&��Q�>])�%�T���k�ҵ�ާ�/��aS�3�P�>�b�DN�]�	)	"4�+��1��"������D^�Nc�LJ��M*cᰪ��C���w�Y���N1P<�(��}��8-���m��cw��m��S�pf�Vw�L/Jc�|�V���ye@��)�4{�밢C#�.\Q���=$�]��|�9gu�G�����&�&y�Q�D���Q���A��C���lW�^߱���7�ë.N�lo�<���-n�;�{����Ng�Ο�L�5�mm/_	�W���^;��!^���=[~A�wV���b�_ŭ��gͱ�;_�r����r���Y�乁}�m�mz|��23&����E�^�������TC��ˑ�H�z�u��dv
/�\L��p�ܶ�}�O����+.t�O˴K�w�޲�T	s�o�PM� �ts+b-�;z�X>B`�0/MK��r��&���&��8jpC���2�s����"��D]�/Zr>�.���9�g��G"�YD0pϾč�e7���>.E�u���З�=�c��.�=m�)�a"�]���7R�˘ ���Y�9��>a5�|47��>>��erH����6�89pɬ^$,����{쁷��	��U���-���ywP�%w���ߥt�{���Ϫ��Ĕ���!�8"�:�u�����&� {������D#����(�I���u������B2*Z?��Hh�V�6y�_)���쯲=�P!\/
��Z��Ӷ��{-��ˡ���h)�$���6lh�oI��O|6o�͟j��������^�t<�]U Z��̐�}�뷏)�(�fP�p�]�(����<=���
 a��0�j�lX/�&,����=4�/a�^�X�p.�#��x�B�]1��n#m� 县�&�,\�.'
�rmEb�c�F%}rx�������1r�M��A&�?H��^��$=X�+G/4!y���廛��|G��7]�ʸ�d�(� �DV��X�^ޔ:O�N#,��� �H���C���m^[��`�Y��S������a��h��tqϑ~)#�^���Uͥ4�~�&�8����SDf�b�ع-?\)��/��~��!��
��^�����+µ�)�2�Шw���a������"�l�����{�Wz$X09��7�!cK�c/���k�q�j\�W�D��E�P�Y�^?�����D�oq�D����NƱ I�D$M'���I���� �M��E���RbvWnt(Zb�_&ц����8l��֕�̅
�D�	a͒`��U.6LT<���L�ľiz4�����0�.!�&7N��p��4F�q�0w>֟�����G[�����rJKk�6MXzAƐ���/������- 3vN'M��@�'��7��q����Ϡ�Nѝ���n����@�_�7{��խ�aL���v����^�h��e�\,�h��r���x�>*�|��&(��Wqe'��,f����!�*�8aj��xh��Uig� ��>,(��w�B��8���M� ��6�Β�v�M��vO&:ßw��1�v�"3�h)4�kN�U�������۵��3~
wX6�\m�0::�Xl�n,O�\,̓'���Eֵw� ��\��7�qfR~mx���y�0�u昉5�h�)�@D��:qm��-ٰ�Swg�����ߋ�o��fV��������eu��2���f޶:0�B0?�I{#�n���N�7
}չ�ϡ̭��V�}\P��u�S7 �OS�����Me!`T�AQ�R����Z("E���S��'v��i��\lM\� #��"`<ǌ5r/��kL^�?�.:�V�����c� �^�&�����0'-6,+�߱���"驡�L��L��x/��e]���o�ߣ_ψ�=���d�\lyW�M�xD��Ȑ�Ј�C�ӯS=N��.�C��x/lS_v ��7Z�"����	��Gr��o}в�����v�<���uI�`\�r�9dm�CcN��
Z~���̆9{��-Q���ɖ����ʦNXo�v$	��5����8̐�~�������}��2��r�,PC$�#����B"+��_�a�c5	��ǹ��	�ڱh�I�� �����)���t�-4l�&&�5jz��$�>G���H#�W#�n���Zԟ{�}j	�����@�6�\�y�B�8<Y�dav�li\1�p(��g�JYh�{����p?~T���B2��D��'�����z����57.ȇ���WE�6�E������6	��a�Y=���k����T�^%�5z���q�*ܼ"噍��Tdhxq�t��v���'c����	�����E�ZV�t�>�7�p�$�˘���W;�<�����8�!t��H��r�g(4�j���b�����uy����F�N�4P�:/h�
L�6�f�j
Y�'�&��/��ku������O��8a��5��3 x�u��/���+��mE�n�7��R�1�jK�4Q�mO�.A����agM�XI˫��hEZ)&u�0G��~o���Ղp0#\D�*:˞�{�r7$ldz�46='a�)�.$����E�>]�FyY��xCa���qF\����f:�(}���ߏ#�-�����w�S��%�e`}Թ�9���9m��k�Sdi�^�n��Í�#���N����'b�Jc�/����h_��S��	�]S+{�o����m��P'Z2|\�5ĂݢK��#S�qh#J�٠���}��D��J��q�U��5��j���i;dV��Q_)IY���gx��3;�����T?_�'�*D�ZA�D�U�_P�U*�g���_��/�j;R�,�Q�/���-��BP2*1{"�nH8�+���p�L/�T�i6�̝����X� ����E��Ct�I�ma�6�����[cIø���z��\���us�^Jҁ���MjkC��(0��ɱ[�7t��]�w�3�U�r�)�3�^��f�+ړ���Te9���i���\���I�=�(�'�O*
�E ~=K��Ω����ؙ@_4?q����NC�?��U .��8d�4��C�W�>u|2�iR��G�^�l�-&YI���Jl�0��Q���ܿ{X%s����&=�.�(q�%Qm��[L�M���H��^m���
��5�/�
�j􂪔�,.�E	���

w�r%}�;V3�.��J-�۲ x�=�&�ќ8%Ov���'Be���,z{����8���r���S/�P_Dq�TԖ�=F
7(*�.>ϛ�����R4��.���ڪ���	�d��)�
G㞰9����F,�cR�â�N���i� cI#�1�П~��Q���_�)3�T�Ŝ*��Oj?�e�~
F{�;"ٓ�L������j�,�����*����n��r}�3Yʰ�J���]|���o.�l爇��� �O���9��)(ޡ�� F���&z2��W�Y�Ga�ǽ�B��Y�?�ް�r|��=<P'V����+�����߰o��|r�min��+Bf����vu��lym���Zx�3��RGw�F�͑Wո\��^����2�=C%��Y�����0�hcc��v&8{o�]�:�/��5c<;�V�M;���{˟�_�1�p�.�2`��9jv����Yi�9P�o4I�U{�����ݣ��T����<F���'}>��?�se~��|
���"�A���E�ʑw��1p�њѓ���3V�/�!@R��IX�`^�2!��y=m�k̿����~�^��ԉ��%��2?��} ?�zs=JY�L�����W>���oY�"�	�G^�Z=O�eAu ��ߒ61��׆��/�{��c�ֱ왐��f������Q�3}6D���u�m��w��r4w0~��D�0��@����P[�b|'.($�7��Q�˟���E`���GJ*c�eI�2��)�#������s<50��[���Y�s���\2�E�Dk����΄�`֛
�C���b��VT�8�Fv�-~����x�Y]�zе�q�z�j��&s�N�Lw�p�ܞ>��B��e!�����W���\Ϻ�g�����R p,����:��Z��H�V�B�.��?(>��Ő7�M������T�9̔��θ��8EiY5��M��~��4L�B�ɒc\�w�zU[��L�,݁@H�D���H��t�3��%��⹡`�4M5t3I9i3�OH��&,��CUL"J�&>��J5纐�Oo�$�qD�
 �"ׂs)��9��	��<	�xn�~h�Xn;��ˊ�w�6iM	'h-��V�S,FkĨ���N�����^�|A[�6d��O�( �-��m���	l�X�dtn�'w�ZYlSG2��X���:q	;��j:|�K1')�7���"�K��'Hg��D����]8��y����e�T���KP�	���W��a���Z�x��r�{�ű���ĵ��@���+Z-�}
zqSe��Y�t���1���i���H�7�A����Sl,�#B�����qD	�sp"cҤ8�D����5Y���2{Y4;��⩮3|OLݵ뼱3��ڧ|h�୆�h�����=d��?ij��?(�E�5)n�-�tj:�g��M�Y"B�����#������t-���f�xDX��F�g�a�}�@]8���9���8k��އm��gQ
|'Ri	n� Rv"=xC3 ����D+��;�˭�
��?-4�5ʜd��1��Y�Y�7?���U�Of
B�\���3�K;u�[�e�߀�=�4 {��ǻGnh���f,
�yM�ͪ����F�H%�k62j�ح
�Z�j�#��^����%!�o�b�,�T����P"@�͙��*6���<�@_��)|�N�{nm���He��ҍg����5F�+��z�wo���U!�
�<q*�ڦ��\��x(̡|&�?�,7�t�;=a!º����-����8�H����԰u��(�P�+<��=Ւ�J㽥���_8r���̱V���3&�׼7��V�V�$�`���R�R��[�o�MG6m�U���Jf��w�1�L[�M"������ԃ	o���Ι� �V�샨%�Ub1��ێ� wl��荃
���M�2���{97+�.!���\*1�^�l���OXcFxarǱ�+u�gA~1rtxo4���p���g]v��cǰ������]lg"�O��~�@؜��rR���f�95 ���F���4��g�u��d�#��* A�+�=V�P6���8��1
9�6��m�f�/��=�=��n��h�af��@ʇ�,���L�k�e���g�'ub��H�Ӡ�W���к4d���h�9�h�J'ICr>�ďr�k�M�>X�rW�?iw����T4.S����Fԍ2���1��0b]0Ѹ�N�n����Вm0�k�A$���M����Q���8��Uޗ	y^�C;�PS;l=���T�7G���{�:�U�X|>����u@��%��\D�?�����p�i��d��T�WǑ��zw`�:gP��&�#e�3�� ��:}k���vg#C�oF7>��p7���
/���� �u�!,խOlA���/K!2��N�A���I4�׶�U���EҞ����cM9�ڮ}�����ɜ��:��H�RՇ��-1xjvj�W3��l�<��	z��hֶ0�g��8�o�V�,B5uWLP�D�N8�F0�h�O�Jk�Jl�X�v�t����e}�B�S�\BM�y�Ƿf�T�}	�%�����|��ػBy�u��dP˱�Rl�G��nq����T�Nͭ˿�А
]��G�t�kc[�����:�q`��ř���C1�^}w��E�@�w����>Y�E!���	F\���wNY�{�:��W��?艺�%����r=4��� �-�M��HԠi�A���)(S?J�~X�pk���<����_d]$'��?8�c�4
���ŝ��OE�C��	��}�I$;�HĮ((�ҁy)�ߤL�d�m�W�_o�{����:���MC��ڨ_�CS9���O͙(��d�8���0kF�����5�u��/�����J_I��7�`��d1%�(�h�`A�oU� +VB@D� �вd��K�b�} �}�<OS�8'�������"Ez�2����1����rs�2spH:`	��!���d�<��R��BR~�l�
V���<�s�ߋ��)��Q?x�9F>�W��޸��o��a��&$�J���}�H�ZgLM��L�pd��y(���H-�����ӛ�h��_t�M��u8W�dc��s �U�X�N�)��^p�i�0�r��&�8#-N�g�y���t�ao�j#aҪ�_�0a���ԇG�?��v���@>��]1������AR"�CkS�s��Gm?d��Sb�B|X� #5 le+��M�y�NP���}��H�����?9~ ����*�����a$7��1>�H~�����8�RF�F���#������a�+���:k�o`�Ʌ�Y����<m�@�L�*f~5�l�8�I$Ҏ,��A޽��T���],g�i���(�]M�1و�=Iz%��&�z����wtDj���t2�z�)�h��q����w7�-S��d;�i���ǖ_��o4��%��VZ1V��-#�5�K�{��i_�^�0�2ԓ���#V��ľ)�BV��eT '�}�#��g���{<�B.2tml{��h�ˤ�!t�O"��5�p"��<C6���Ԧ�z �EQ)>�}�#)b�wk�m��L'3�]:%��uo�{�l�����eQz�p;	�AZ}˳	L^��N���q!�;g�b�>�*5����7V�H}ֆ.�뙇�'��0�ZY����-랂�\;�-Gf�g�A�"Gg/R1�'7�MC�W��M�x~��������L��M�FH �_�X�u�	V{L��� (�L���IDW�&�{k[ځ�P*H���f#��^�.l�DINu/^���B�Suo���f��y�)p��`O�n�v4�4���'��E���{���n82z%����c:;�A
j�?��69�}����ؽ��m�TR������h�ݰdB�b~RE�ў���^�nt��AH.j��<BP�`L@�+7���E7�Ğf5��u�Ƭ�N�[�:^ק�E����lz�m>-��Eʎ�5v�'vSc�@��pl�$G���`���H"#(!=�׬�r���m��M
HOD--wq�S��V�lٺ��=9�'�+���q|V�jyk>`�n���~��SH�1m'�_5&��=����C�S�z��ŀ��.���I�P��;c�8>o�+ޗ0w�"M�ߏ��z��f�}�_�����5v��,�{Ȗ ��T��kl��-�uOĬ��Sr2˨�f|~HHN�t���ɮ���I�8�f5�	h�55�_�:��C��H���-���$4�D����Qt�����D���*�g�]�0mG�34Sp<��R�]a���?}Xf��K�F�V�<$c��w��SI�(���>-I��^	�=���0&<���&9�DK�ܽ��rO �&(DJ�9��_]�>� �GC[ք(�8D:s�2�!f����#������s�/)7C�,Q�8+�p�>aRv��屨��N�?��M����iU�n�?EM�P���O�,y�G�F�!��g=>���?��^��Ǻn��^�'�~z�b����������>&�WB�YB;lz6�(d���)���o�-�3�D�x�����:�7P����\m�Q�0��V��f�qk^;;{%9�!�{g��ב������T�^�뀈�z��AQ�A#\�v���eD�4�*�i�
~xeK�>�I�s�&1ܰ��� h�ou>r�:�,�C.f;#�0���T���	B�P�3:m�g|��I�I���jo�7���&n����хz|j�����8.,B���Q�ez����o�����l��f 53`�� c��0�~�^r�O�R�5 rXJY0�8�i�j�IQ��nI�
�*2��*;\Rhs7 ��BA�Hі3:V��hynE½RP����^��:g��9��*��	�����������8S�_�|��t�t3�aP.	���!�Ln\[�ʁD�x�Ò]fi`�q������,c_T`T�3�v�m�k���%������|�x�!p?Z$�v�I��/T���F_��ay瓫n]��-v�R���;��,�����`�\<lkߑm���?3�ݾ���7�6�f�����AwV��D�nr$�]�B�	�!N4��.�l�U��XWd�d�9L7��%��z��n_���]��Ŭ9�����6Di���T�IAG�+
c���pk�2\�TzGDm+�>��V[���$6��>P�,�K��R�sʸ�/�̹�G.â�U�@��)����)|�M�Ҡ(��wU%���77V����x��]�Y]]J1@xF�v�����:K���q�CB��/X�zd���Qw�У���%5��\�MXg��
�������`iʩ���U��t� ���@�pY�-1�N�f��R��֊��d��c���F�>>!���/c@�QJR���+R�׺���4aK�6̩���Z�UyG�G��˄���Y������#.:Ǵ�\�x��A�.l;q()ˤ��Z[�{J���7b;�9r��]���e��R�:^A��:��S��7O�����`ф
c�g5��ߚ�h�	��E;%-l�$s��5��X��y�g����FȊBy�xnڦe?��V1S����wU�h�A�����f��0�d	�����N�ꢁ]t�:�Rd�P�|C��nP0����EF��E)�t��c^���<�q������i<��J��0�(ŋ����9�\�B�o�܃�8�WPs�JZ+kQq�$�=�oU�"$�o8�:,C���l���H�w��`W9������4�ѳ�'��!oO*�v��)�󮉡i#�}<�Q���	�/�ӭ��L�s�2.W �"0�'9���J�x��n.�i����Nx�,���g�	�%<��3�_ �M@D�D�F�{>�8��e�f�b�� �S��5��EH ��9(0���̦qSz�ǐ�j2���첻� $f!n��~�%x�K$�%3�#�`�
��;�ҡ�y�%�%,5�`,Cv VK�G���r~s��`�/��u�<ԧ���侕-�������ӫ�t�՚^�S;9z�xto�Z:ڲ| ��r̟'���]2�ԒĀ�\�ܯ����T��ux�6F�>��Z%���H`1�d#�����I�+W���f�(7�����]�kW�ga���j��_��-T�v�6��z����i`�I?7����Nj��y0�{
m���z�j���P�eR��FdI�ɢ�nf|)X�v�P{��~KD0�t]/Ƚ=9��Տ9m�ô�EJ��@�I�@'4@��U��]�;�$��bJu8�����9��v�����0���7Sa��� �i� �H1�c��55_3M3!� l�I��:D��>��dHp{�P:�q�DV4W��M!�Иt�nĂ��=�7��-�6)7���m4w�<0��M�}�?#�g-�]���D��.��a�]��x ����g�*�*XZs��(�l}HV���E�&v��z��Q���C69a�?Af@�)�j��0�����=�QPGl����$���Th^���(P�m�^�C�H��ws�n.4t�0�7<�àv��VZ�Q�hX��*ڸײz�����[h�P�N& y�S-�~��c�����V��~)B��ɓ���6R�!���яR겠�-a�M��zy�u�u��`}OS�ٗn�b55Tn{)ۡa��t5����"u%Fx�,B�4n嬼��no]�A=������NN�*��<�15�K�)��������V9�"F�(Q O�#��9ܱl��?������ �֧
�>}"Y�Kn��0�[�GV�cg����X8���?V����)��e0���r�G���5J�l/S���%�"(d������L]���(��WnE�c� c���[�2%8�C���ߩ��|�U��9�A�����9�0/�=�I��D�A��R�;�v�t�� 􀔶/�R�gy��߫g��E.�d^m�����{Y�T����%�_��-j��
v��x�I|8b_��d}���X�� lY%��9�n�([���h��c����-=�|�4 �K� ��3�>��T�Q	��:�����
�r��"���U�u�+st��}���P�=׉���ʽhOǏ�K1?��z5����!$
�h��&d>�p�qQ�_\��#�{u.p���`��3V]��#9$Y���AyUi�Y1&[~�e��rZf?M&B`��<�����;��]��q����9���*��c���[o����q��T䎌�Q*��1��	�7/���F��p�[��	p�d��wd�ŊE����=I���u�X��;��������i����=��f�Ec��}_8a� |�+9���G�J�#�cɥ�����w�5�/#�P�5�8��/��VJ�D����^b�@�9OAć�9e
X�;|kiב��w�'9կ7 H���@޹A)`�C-��T�4����'R��J<-���c˜��	a�5x�&��G�YV(�&o͑�5_Z�lԥ}�S��,�����	�+�^�SN�BX1�>�$qt��ģ!�5��%
Hר*T~��.�F�&B��D�Ȋ��H�KSF��:��>��4s�_��;�cT�x�u�91���8``�D�����_$̫���RbK��g��6�G�N�d'���^���Q+qz�t(zZ�&\��Р�2p�;Ep%6r`�U��f "6���%,�xx�u坈2����іk� lWP�����/$����5������o�+��!�SP7�����՝=�<�z�c��K����i<���_I!���u�v;8�>� �jv�o��ƾr���B����W��~=�	��+*:c��@��,ў]G
A�鳵���n��#C][Tw���*[�������?�n2t S�j����T�J��~}y��K�5\�ښ�-��!���%��;�T�(�blZ���L��ǹ�@����LP)��G�p��EC�����gDC�3@VF,>��s�Ǵ.@P&�g�R ���X՟�Y�7ml��ϵȧ)�c�;+������~z>8���ڻ����B=�u�i�лC���С�xS�gFD®G�o3;���Xe9��;�\�>���	�6!@��އS�(��_t�xi��Pj{@{x��N'�!5�ux��ti1V@d��7J�r�u�]Aw��9��ܵ�5���c�u��9�C}w�� o�i�\ �e	C����W%�2̪|��
d�l���|65��v��q��&�\9�a�b:\|x3�_���m&~��h�`��
^���� Q�Eg��|�ٱ��x]�I�t1�jk
ړ���hxd]Od��Q5@��&>K}�K����Dh OD~G��q\�Zޞe�>��"�������0G�Td[(6}�"�Yw�3%ґ~�ud���Z��G�o���y`h��-��{2/��r�V�؟�Usa4G�X�l�S�B�xA���g-�O��>��ph˞5Sr&����b��a�i-ߚ��`Q@��k���p�drJi_�p�ڙ��r�gA��;�{{�YVKp�ѐ`W���Q܅�\)��R�Ao�)�~ij���OV��{!?Ӭ�6������T7��V]�)�6�(������(��j� 4}�.���&94��������SO`�ЉBi�Ϭ�h:��J�ӌ�s���������%�����k����̇��Yi�O�֦��
��rۗ-,�D�F6�T��g���4P]%���]j`=�\��U�)�����x�S�^�R�
ؕ�V�=����g��+R!�ؚ��mD�|�¸B,���	K�����5R����#�����.c����eľY��;�<�k�S]2�+�Ԩ+����v��؜�W�]�8u\0	���+o���a�+�l�vs.�G�H#����@�L��>�Y�����D����h��ǁ�!�ݿ�e�J������w7�\�#�Ű���<?�R�j@X�*�T*��"��;&r��Y@���f�G���&"M#'�x��ϊ�3O�D�����(��=��J��T2�>@wЀ{��*ըb}Y�� �2��ї���o�"8��1#؅�
�����%�geL�P���2���"\��^iO�DML��՝R(V;xd�k(k�-v�o��Yo����X2^Nth����E'`h�	�s�
6(B��7��h��S�<H�To�-���q$�
�1Z��e,:	AJ��
����NEN7�%P�tO4�l�|�����p	����,�z�i��w8��hHk��M����b)�����{Q�>A��N���w�4'Q�ßP����~������k��g~����H��ߟ�g�&��Ȼt6u�=��',~�>�a%�:�4�N�����M�r;|���2�=��O& ���H��I�6���u�|h�(�p>��-U��F���ž�G�W�=��E�A�Gd��l�_)�j&#ݫ�|s#+J����<�Xi�Z���o�|�;^#�bR��~H=Kt9F"�R����p".�W�%u�E@��!|uW^�\�я����ݙ;��W��nAh�
�e/��p��<�M���Z��W�T����Vm��!a�8\9��B��>�@b��Թ�~���j����?��H�`]:�f*�2V�ܷ�2U��
��ZC��O�V.�Au^P�An�/�XD�Ɓ�������Z%����!͒"S!����m/���g3=�Dg��B�HU��c�x���*��{�Њ,�nl	�8E�̝~���W+w	ɮ*U��OQ���=�w�Vֳs��Y���+$αO��]��0�o��Jvg �`Cp�r����v���\��NK�n8f�2�^x�6�8����ϙ��6�6L�<p��� ��	f7��Ĝl�����ƃ�Ge�"rBxX>��n�[���It־˲����.���Ї��V���uXǩfy63abG��H����N��������^���{�D����M�ձ�kCwfK��6	�`' �a���<*Y��� �"u��,��Y�u
v���'����� ��kf-[�{W8u �6ou@':xS��D�
�tL:����D��v~Y\�P��a��n�: ��`�W U�w��.��v]׈Ǽ?Sah	�Wa��-{;W���*�ǃkc�D�w5`�0�>
UW��X��nq"��m |��W�M����d����7����K/X5�q���N�[��{a��jP�ʞ+A:�r���{�g~P^���ٚ�g��p:5��iàc��-6�dy�X�"1�Q{	
���V=L���JKs��N�ZF��;��=#��֥k�-��A Zj��H!O�z'��#���`�P?4���$�Id�}�� W$B��{%׏@����d�y@�_ �V�)ξh���b{�ާ�W��kv0>�^>�ZY���<��s�'s8�9d�1��4�.���+���6�|�>y�E&q<aܖ"J����oꃵ;��R�()�ݭ����/�����P�=k�X^���˦Qw.���L����K�I���f��8Et�3�/�P�&��vڭժ�b.���	����}�_�؄2���Lκ����V�,�HyIU������
rt��/[�<���"��N������R��F�o�o�>Q6E�g�Jd�\]��Y�����ǅ��[B�N��#|xL4"Ɂ��
��M��|t���އ���^��M-V�P��Ve����َ�2�h�����i(v�J�i�Y?�lk��3V�����,� �K�0�
L=�s�[���Ui:������¯C~�f�M�I��z䳶��rC$�,B�P����4ěf�B�6/5�1�B�H䴉�\�]����u��HD8�y�4njN�*� �h����4����?Zˎ�F�p�}��;��!H1�iM��� �5��n�'��~k��&�b	����l�NӉ� ��?5a	62�&����`6P��㺀���&n�|����3E�DL��!�g�(�S���|> ���˕�qC��+uǙbe47U�)A�V1�Q�/:��1���h6�J�2�`��%W�R0H�F��)�G�� ��ޣ�Z��yZ����)7b�n�ޯ���W� �|/�:;,B4�6����ǻ�ҨC�Ք�Y�I�t��_�\�����ʲ��ۚKf�U��俛��E������_�6-��D�I��W�>�}�ds�+�m���~;r����4��N�.��|��l |�ʥO~���C����ȟ|(�*��)%!n����W� ��)�uR,��!�??���S�^1�����"nU.yAS�ˉ:$sZ�Ǆ �`�]KF�`HN	�}�Tni��hӴt2�ba�u��6Ƿ	aA����r#���|�q�ˊۀ6�ʍ� ��:nl%+n��)���ً���W�Q%�z)�,��8�E4<D���W\H�:�Ǉ�{wd�B����Kj�,�ĭ9�(�Es@@n��T/��
RƷ1 &�A�|͐��	{��lw�w�E�Q�\�u�y���u��B�.�J�0JA�*�W���Q���6�W���qw�+&]LS�Fв(�J�V\�������+l����<ڀN�\�t�ƧO�-|%O��9�g\�U���:��6��D�T�s?U���aHr�����D�OIo�i�Q��#�����9>ZR�~m�J4h��o��'× kX�=9�8*�Q�E�T��ˣq,�o�+��`�XP`���L��kE�స3�J �Ruˆ��� Hc�J�S|K���j�	�_UT�sW9�5D��,�WK*ґօ|P�y�N�ុ�K�F� :�g�k[�Y];AG& �uG���{t:��͜U0�$�N��$������� -i v	輘-FK�\�竭���Gf������f�pzg�@������9��Zm�i�s}���Lo���!��n�i��^�\�@�+�ȧ)�j��/1K���v亢�,�"?�������.�G?�b�c�� K�!;�R�D28	��Ua�2�/BE� ٳN�j����6%�[�u7�C��ՊU��1*��I�?�lkp���q���5�c쐶�gb%so�����$F��f&�[�[���0�b���^���ϭ:L��ny�[K�t�9�D��H���=��Yⵚ�$}BI��l���ك��}��"n`Lʙr	�&�k�ԝ��N��&vz"�2��@�q뭱��}+�#m!.D�X� 
����b���8@�vPU����,�F���^MMN����Ind�6�>a���&�d�/�i�@sL�7��>��\���d/���ӛ�qE�J��Whu�z���nS3#��}d������d�tw,��t�L6]�����}�>��"Z�C�G�8��Nc�J-";{�:-pp�V�҂�� �Dײ�����2��{@��U�:BD<i��J_�mδ��ې�f3���l��!�l�{���Ml,��X3��]W�$녥����6�,GN��M����*6sǠ�9W) ����j�O>|l���WX�/#pqm����5j��t�zZR%F��J�˪�Z���bj���$ M���[�v�mB�|h�]f�O�����6N�p�Ъ0}ۜ_K��6����2��2�z�	R\�ʼ;�$���TMe�r�A��w4�����H���܂�iD%�{�7�2SCF��:Ǒ���U���:~�v�%�I���WH,�S�\iBx��L/]?=Z�c��S1�',�6�o�ɩ�q'9���9�u�¢�����>��M�{���;B,Nq��a_ �l� �g������ۄy�3a�O�M�R���m�3^:����[�=劜}j��Yʺ� �|��x�;W ��rY�%������PhF��E{�sa���6�����}�(Ki��;\�Ll�9�.�}�#�|���&i������d:�M�o9�x�T�5g�&\��R�P;z	�oD��"��{
��&��������v��o�5�Z�A0�q�sO�N�Q�53��V�Q��h9�S���d�z���b踱KH���r[Ts\/�C���Eu_���s#����n�hLj+/o��!�bhT�+��#�<�wx��8��nm��U
�i��|��85o�,8J��+5]��=��;U��yo�l����?�@��}��K[O�0Bx�t�>Bb�G��&y�)]ҭ��ܔ�	x��YG�R]�i���*w�{58T�2ꬋFE^�/r�ԫ�����17�Z��vR�j��ӟ��˂/R���^�H;0�B �����Ll�>�?_��$w[p��v��*t��H�� %�a������9.<�C�krl{�����V*S�k�>X����~=���m�?�fj	kg���~�aLlF��B���Ug�f��ӏ9 2˺�����2S
� ��c���磴���n-��FA���/ 8X]�|;����݉��>Û�Ⅲ������J�k���X�T����_O W��߈UGJ��M�H��/:���9��C�X#zK��Kk�P��C�����}�V������&���i]ir�,L����M8���N�I_�~j���h],JX$�b�w0�P�dȢ@�^+7I�x���\�e�l#j����=A�R.0)[J�=9�P�Pն��k./�K�f`�a�?�TWh�O��]��l��#C>o')�x�	���ȩ`:����ߚ�'S���0U[z�p^�Q�:�iF�_�Aٳ�E��������+��P�' y��8�(z�����<�ٗ��fj$� �^y��r�i����G�0ak�_�����
q>�(��ȡ��=����I��֯����6����o+`��J� �1�^D�>"����X��z��@���Fy3B#C��A��i��wA>��'��o�=}�r�\�l����a�H.�G?�r��%�a���X�%J��Pe!'vJ'�W���S��@�{��ڸˁ-�d sz��{��"E�Oy�0.i� � ���Œ��N�!ї�D~��l�����_N��� �T�KfA��9<������0���zdR��X;�5	׿�Iޥ7,�^��.x:�x�#_������$���٧ǞX�w¡���Vhږ�%1b�13 �P����#�@ry�� �
���Y7�)��O�(��e	ס�!E:��>�ˀSN�r��7��U�'��c�/�f�?j[�rg�}pY�M<q��G��BW�5�Hv �@m�(4�V�'��4Y��{��2^��3��.��z:i��q>�,f��^�M�N��`���QU:���\Ў:�:J�,Nn��K|��ĠcE���ɦx>'f~��!�T⥅�c��]� ��j��1Nv����f�Lng� %��eW���ʷ�2?$��zxL���%�xF�/x�?���q|O&l�h_�E�J��J�b- � ���#�K(|���CU�G�Ջl`�M�ag�/(���EK�odf�+�����8��������48�Y�
�swz�� �v����F�\�d��^*��\�]] �R�l�R'����w<�����j�t;c�|������O6r��@��|�tݘ%8��Z��zQ%Pn��?5o4�#��a�ԏ�NIP~M?��k��v��i�rx%������~l^��; 
E��
�ز\���J�'V<��� ��؜z{�3@��\����Fs�ESC6���*kD�uOM[�?<�#����9
��IW�9�!�z�5A8�\�s��@}X��F
F"-^��$�_.䔑'�<�(7�������(4_��5��	����4Aʞq=�>��ܸ���*&	%��ۣ;�=��G�O��@�� ����J�X�+xUYxEb��. ��vٻY�F�2a��,����5|��4Z�CL)$ž&�}R�`�Ҥ�d;K=�st
q����3������iށ�U��*Y�n����^��b Eep�;(�ɘ�g܅��Ĺ<j�ka[�'U�_���֨uj�Z(7Q�xT\�>2~�4Sz۱�Ԧ=���>���w�!��i�g���-����X@3��
���;Fx@1����R�����?\WP-zK3�G���<�i��򫉘X������e�QU��p��x������mX�����(\|-Bj�@�ҋ�Ϯ?KǗ�j��z�P�7��E��Q��L�����|��߭� W���!v|nt���Z{iYwBީ�p">�R8��������m�ĻbSN�7�Et���:�#?�~ X�#ɠ�h䊜tU��&s2�9g虻��͊�����������45)���^���Hk:L����VU����ϡ;���s1��@��S��ѯ�{E���`��/��A,7��f��K!��W�y<�t��L�� wgGe����<��u�xW�� �N��:�o�y���x&�1�Z1��``����^^6ώ�p ��~�p������n"L6)�\BN�xU<k�7��H4��?��{u[%n����逋�����	�驅h�PT)����^f&�\�C+��So�'�r���%Ђi��DJ�l��v�=ȃ��X��%Nz�o t�P)D����ֹ?������PY6��;C�GVN(@���b]���� 	K�`'�P������%~�b(>g*u^�������rv+?�E`��N;�b�,��e�<9�Pާ ���|'-y�N���ؚ� (=�9,�*ڡ�-$� �N��Q��?�� ���wm��d��C�%�A���,]y�>�l��+�R�~�,�1�/���Q�w>e�R."$�Jb��&�Gu�[;���J��e�Q�\�K��B� ���	Yx�h:&�c�b�4h!���X�M���@<�y��u�,���C7h���b��!�mD�5x!�}�K��2G�պx�����wRpf($��� .Fl��42���[P�B�w�-eG�S;A�bh���O�kE�Q��¯V��mu�=����,;J��	G��L��.玔�L@ yJ��OF�����\��/I�<�C�TE�!�2��gQ�� \���#��\]s���z�@<)��JU�L�~Xf^Ȝ��M��SM�ͦ��O�aaU��%�C~�!S����/:�)3���1���ϧ��a�P��S��h3�l�?�\xr�n�U����lZ��_�0�}�����Isyuɱ_ �2���3�[�5���2+_�i������R�1,q{E��ω�z(y޶�;Hua��EYA��w:PN�����o��������vhm��@?pe���tj����V+	w���)J�<�Hn|��Ġ!�0�g?тu`���l�Ϧ�ĺrx!�����1����S%��"V�!��ţ��F��jv�pM=�V�mJ������t�ߔ��OZ��EeM_�48%��Y��D,B��@e��#�[cp��k1�~:����r�/��i�5;��g��O���_����`�<I��=&�X��w��e���R�@��*���!�Ӳ�������D������2��ί _���n���3�!���(=�h�.6��n�UVh�j�Rb�M�.�2��ٸ��%�X�9��')� ��	���e=0�6�lyTd��
N�#G�m���K�6.w�Mq:ɧ.�=D� ���$P�Y)Y)�#/���>d5-����<XM���4�~���,s��K��5c��=�́_�]��0lj~g�́OXǩO�"r�,����:K�eBl���"A�'�ׄ㦋��Qr'mכ? :��� ���X��7IG&=��K+�ۚ�b�dW[?���?h���AEsC�?,��v�O�����������wŦ��k���q�h��������n���u�J�=��S7bEոf=6���q������jUI�}�i���a˖6�O�3��~{d�h�WJ��%���Kl+�^������]�"gUm�˚����.��(p{F+�3O譨���*�wqPquE�Y/�Q;�ĊH�]l���g��r�ҕ����ik�]<7m���%ꕿ��]an�G�@�^���<��V�!��
�ؑpe��r^c����ҳ���!F{u����q��R�>�7�+��O���
�R}�pS K�O(��:}���MB�Y��e m:^�K�#(4�7�s/������P�&�#㧤��bttj����P)��hp�m���r������d�o�%�垲�m9\��+'��Cu����_��#�ɖ�V4.�'!��0"��e��d^�Yb�:���Mw����g3�i��m;�,�W�`�x����K&�N�)�*K[�朚� ��缟��Ӌ��$0w)q@��5��m�~'��06����0�#��9ʰ��Q��h�&BW_��O�~"`e$��Y�e�42a�2�*����3�F] ��"Fm`�Pv���J�\�+k�г���m��.,�k4��_S�������ƲDQ��]���/1����e,�b�L�E����2�k��@�^~I|�ہ���!��z���2K'�$�o�����u��%L��~�}�פ����K�ʯ��Z7x�jW܍�ȅ�9*�*]˞��N�4)Ӳ�_�p����`�C�T��B=$]�V6�����$���U���\�n��VI��_�<�&	�G��@{ *�G��y�c���S��QwG%����\��T���